library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tempest_cpu is
port (
	clk  : in  std_logic;
   clk_en : in  boolean;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tempest_cpu is
	type rom is array(0 to  28671) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"02",X"BB",X"5A",X"30",X"50",X"EE",X"3D",X"A8",X"4D",X"20",X"C5",X"92",X"20",X"34",X"92",X"20",
		X"2B",X"90",X"20",X"31",X"A8",X"A9",X"FA",X"85",X"5B",X"A9",X"00",X"8D",X"06",X"01",X"85",X"5F",
		X"A9",X"00",X"85",X"01",X"60",X"20",X"1B",X"92",X"20",X"C5",X"92",X"20",X"8F",X"92",X"20",X"6F",
		X"92",X"20",X"46",X"92",X"20",X"9F",X"92",X"20",X"AD",X"92",X"20",X"6E",X"C1",X"A9",X"FF",X"8D",
		X"24",X"01",X"8D",X"48",X"01",X"A9",X"00",X"8D",X"23",X"01",X"60",X"A9",X"10",X"8D",X"02",X"02",
		X"A9",X"00",X"85",X"29",X"85",X"2B",X"AD",X"21",X"01",X"85",X"2A",X"10",X"02",X"C6",X"2B",X"A2",
		X"01",X"A5",X"2A",X"0A",X"66",X"2A",X"66",X"29",X"CA",X"10",X"F6",X"A5",X"29",X"18",X"6D",X"22",
		X"01",X"8D",X"22",X"01",X"A5",X"2A",X"65",X"68",X"85",X"68",X"A5",X"2B",X"65",X"69",X"85",X"69",
		X"A5",X"5F",X"18",X"69",X"18",X"85",X"5F",X"A5",X"5B",X"69",X"00",X"85",X"5B",X"C9",X"FC",X"90",
		X"05",X"A9",X"01",X"8D",X"15",X"01",X"A5",X"5F",X"38",X"E5",X"5D",X"A5",X"5B",X"F0",X"02",X"E9",
		X"FF",X"D0",X"19",X"A5",X"5D",X"85",X"5F",X"A9",X"FF",X"85",X"5B",X"A9",X"04",X"24",X"05",X"30",
		X"02",X"A9",X"08",X"85",X"00",X"A6",X"3D",X"A9",X"00",X"9D",X"02",X"01",X"A9",X"FF",X"8D",X"14",
		X"01",X"4C",X"49",X"97",X"AD",X"26",X"01",X"A2",X"1C",X"CA",X"DD",X"FE",X"91",X"90",X"FA",X"A0",
		X"04",X"AD",X"6A",X"01",X"29",X"04",X"F0",X"12",X"AD",X"1D",X"07",X"C9",X"30",X"90",X"01",X"C8",
		X"C9",X"50",X"90",X"01",X"C8",X"C9",X"70",X"90",X"01",X"C8",X"A5",X"09",X"29",X"43",X"C9",X"40",
		X"D0",X"02",X"A0",X"1B",X"84",X"29",X"E4",X"29",X"B0",X"02",X"A6",X"29",X"8E",X"27",X"01",X"A5",
		X"05",X"10",X"05",X"A9",X"00",X"8D",X"26",X"01",X"A6",X"3F",X"86",X"3D",X"F0",X"03",X"20",X"B2",
		X"92",X"A9",X"04",X"85",X"7C",X"A9",X"FF",X"85",X"5B",X"A9",X"00",X"8D",X"00",X"02",X"85",X"51",
		X"85",X"7B",X"8D",X"05",X"06",X"A6",X"05",X"10",X"1B",X"A9",X"14",X"8D",X"05",X"06",X"A9",X"FF",
		X"8D",X"11",X"01",X"A9",X"16",X"85",X"00",X"A9",X"08",X"85",X"01",X"A9",X"00",X"85",X"9F",X"20",
		X"96",X"C1",X"A9",X"10",X"85",X"04",X"20",X"AD",X"92",X"CE",X"05",X"06",X"10",X"1B",X"F8",X"A5",
		X"04",X"38",X"E9",X"01",X"85",X"04",X"D8",X"10",X"04",X"A9",X"10",X"85",X"4E",X"C9",X"03",X"D0",
		X"03",X"20",X"FE",X"CC",X"A9",X"14",X"8D",X"05",X"06",X"20",X"AB",X"B0",X"A9",X"18",X"A4",X"04",
		X"C0",X"08",X"B0",X"02",X"A9",X"78",X"25",X"4E",X"F0",X"34",X"A9",X"00",X"85",X"4E",X"AD",X"00",
		X"02",X"A8",X"A6",X"3D",X"9D",X"02",X"01",X"B9",X"FE",X"91",X"24",X"05",X"30",X"09",X"A0",X"01",
		X"84",X"48",X"AD",X"CA",X"60",X"29",X"07",X"95",X"46",X"85",X"9F",X"20",X"96",X"C1",X"20",X"C5",
		X"92",X"20",X"34",X"92",X"20",X"31",X"A8",X"A9",X"02",X"85",X"00",X"20",X"AD",X"92",X"A5",X"4E",
		X"29",X"07",X"85",X"4E",X"60",X"0A",X"AA",X"A9",X"00",X"85",X"29",X"BD",X"C6",X"91",X"85",X"2A",
		X"BD",X"C7",X"91",X"85",X"2B",X"60",X"00",X"00",X"60",X"00",X"60",X"01",X"20",X"03",X"40",X"05",
		X"40",X"07",X"40",X"09",X"40",X"11",X"40",X"13",X"20",X"15",X"00",X"17",X"80",X"18",X"80",X"20",
		X"60",X"22",X"80",X"24",X"60",X"26",X"00",X"30",X"00",X"34",X"20",X"38",X"50",X"41",X"90",X"43",
		X"20",X"47",X"10",X"53",X"10",X"58",X"40",X"62",X"60",X"65",X"60",X"76",X"80",X"89",X"00",X"02",
		X"04",X"06",X"08",X"0A",X"0C",X"0E",X"10",X"13",X"15",X"17",X"19",X"1B",X"1E",X"20",X"23",X"27",
		X"2B",X"2E",X"30",X"33",X"37",X"3B",X"3E",X"40",X"48",X"50",X"FF",X"A9",X"0E",X"8D",X"00",X"02",
		X"A9",X"F0",X"85",X"51",X"A9",X"00",X"8D",X"06",X"01",X"A9",X"0F",X"8D",X"01",X"02",X"A9",X"10",
		X"8D",X"02",X"02",X"60",X"AD",X"5B",X"01",X"8D",X"AB",X"03",X"AD",X"5A",X"01",X"A2",X"0F",X"9D",
		X"AC",X"03",X"CA",X"10",X"FA",X"60",X"A9",X"00",X"A2",X"3F",X"9D",X"43",X"02",X"CA",X"10",X"FA",
		X"AE",X"AB",X"03",X"CA",X"AD",X"CA",X"60",X"29",X"0F",X"9D",X"03",X"02",X"8A",X"0A",X"0A",X"0A",
		X"0A",X"1D",X"03",X"02",X"D0",X"02",X"A9",X"0F",X"9D",X"43",X"02",X"CA",X"10",X"E6",X"60",X"A2",
		X"06",X"A9",X"00",X"9D",X"DF",X"02",X"CA",X"10",X"FA",X"8D",X"08",X"01",X"8D",X"09",X"01",X"8D",
		X"45",X"01",X"8D",X"42",X"01",X"8D",X"44",X"01",X"8D",X"43",X"01",X"8D",X"46",X"01",X"60",X"A9",
		X"00",X"A2",X"0B",X"9D",X"D3",X"02",X"CA",X"10",X"FA",X"8D",X"35",X"01",X"85",X"A6",X"60",X"A2",
		X"07",X"A9",X"00",X"9D",X"0A",X"03",X"CA",X"10",X"FA",X"8D",X"16",X"01",X"60",X"A9",X"00",X"85",
		X"50",X"60",X"A2",X"11",X"BD",X"AA",X"03",X"BC",X"BC",X"03",X"9D",X"BC",X"03",X"98",X"9D",X"AA",
		X"03",X"CA",X"10",X"F0",X"60",X"A5",X"9F",X"C9",X"62",X"90",X"07",X"AD",X"DA",X"60",X"29",X"1F",
		X"09",X"40",X"85",X"2B",X"E6",X"2B",X"A2",X"6F",X"86",X"37",X"A6",X"37",X"BD",X"07",X"96",X"85",
		X"3C",X"BD",X"06",X"96",X"85",X"3B",X"BD",X"05",X"96",X"85",X"2D",X"BD",X"04",X"96",X"85",X"2C",
		X"A9",X"01",X"85",X"38",X"A0",X"00",X"B1",X"2C",X"8D",X"5E",X"01",X"F0",X"1C",X"A5",X"2B",X"C8",
		X"D1",X"2C",X"C8",X"90",X"0E",X"D1",X"2C",X"D0",X"01",X"18",X"B0",X"07",X"C8",X"20",X"77",X"96",
		X"4C",X"19",X"93",X"20",X"83",X"96",X"18",X"90",X"DD",X"A0",X"00",X"91",X"3B",X"A5",X"37",X"38",
		X"E9",X"04",X"85",X"37",X"C9",X"FF",X"D0",X"B2",X"AD",X"6A",X"01",X"29",X"03",X"C9",X"01",X"D0",
		X"1C",X"CE",X"1A",X"01",X"AD",X"60",X"01",X"49",X"FF",X"4A",X"4A",X"4A",X"6D",X"60",X"01",X"8D",
		X"60",X"01",X"A5",X"9F",X"C9",X"11",X"B0",X"02",X"C6",X"B3",X"B8",X"50",X"35",X"C9",X"02",X"D0",
		X"31",X"EE",X"1A",X"01",X"AD",X"1A",X"01",X"C9",X"03",X"90",X"05",X"A9",X"03",X"8D",X"1A",X"01",
		X"AD",X"60",X"01",X"4A",X"4A",X"4A",X"09",X"E0",X"6D",X"60",X"01",X"8D",X"60",X"01",X"AD",X"5B",
		X"01",X"4A",X"4A",X"4A",X"6D",X"5B",X"01",X"8D",X"5B",X"01",X"AD",X"6D",X"01",X"09",X"40",X"8D",
		X"6D",X"01",X"AD",X"63",X"01",X"20",X"E0",X"93",X"8D",X"63",X"01",X"8C",X"68",X"01",X"8E",X"54",
		X"01",X"AD",X"20",X"01",X"20",X"E0",X"93",X"8D",X"20",X"01",X"8C",X"18",X"01",X"86",X"A7",X"AD",
		X"60",X"01",X"20",X"E0",X"93",X"8D",X"60",X"01",X"8D",X"62",X"01",X"8C",X"67",X"01",X"8C",X"65",
		X"01",X"8E",X"51",X"01",X"8E",X"53",X"01",X"8E",X"52",X"01",X"AD",X"60",X"01",X"0A",X"8D",X"64",
		X"01",X"AD",X"65",X"01",X"2A",X"8D",X"69",X"01",X"A9",X"06",X"8D",X"55",X"01",X"A9",X"A0",X"8D",
		X"61",X"01",X"A9",X"FE",X"8D",X"66",X"01",X"A9",X"01",X"8D",X"4A",X"01",X"8D",X"49",X"01",X"60",
		X"A0",X"FF",X"84",X"29",X"0A",X"26",X"29",X"0A",X"26",X"29",X"0A",X"26",X"29",X"A4",X"29",X"48",
		X"98",X"49",X"FF",X"18",X"69",X"0D",X"4A",X"AA",X"68",X"60",X"08",X"01",X"14",X"50",X"FD",X"02",
		X"15",X"40",X"14",X"02",X"41",X"63",X"0A",X"04",X"01",X"09",X"01",X"01",X"01",X"02",X"03",X"02",
		X"02",X"03",X"03",X"02",X"0A",X"40",X"02",X"02",X"41",X"63",X"03",X"08",X"01",X"08",X"D4",X"FB",
		X"04",X"09",X"10",X"AF",X"AC",X"AC",X"AC",X"A8",X"A4",X"A0",X"A0",X"08",X"11",X"19",X"AF",X"FD",
		X"08",X"1A",X"20",X"9D",X"FD",X"08",X"21",X"27",X"94",X"FD",X"08",X"28",X"30",X"92",X"FF",X"08",
		X"31",X"40",X"88",X"FF",X"0C",X"41",X"63",X"60",X"41",X"0A",X"01",X"63",X"C0",X"0A",X"01",X"14",
		X"00",X"0A",X"15",X"20",X"D0",X"0A",X"21",X"30",X"D8",X"0A",X"31",X"63",X"D0",X"02",X"01",X"20",
		X"A0",X"02",X"21",X"40",X"A0",X"02",X"41",X"63",X"C0",X"02",X"01",X"30",X"04",X"02",X"31",X"40",
		X"06",X"02",X"41",X"63",X"08",X"02",X"01",X"20",X"01",X"02",X"21",X"28",X"03",X"02",X"29",X"63",
		X"02",X"02",X"01",X"30",X"01",X"02",X"31",X"63",X"03",X"04",X"01",X"04",X"00",X"00",X"00",X"01",
		X"02",X"05",X"10",X"02",X"02",X"11",X"13",X"00",X"02",X"14",X"20",X"01",X"02",X"23",X"27",X"01",
		X"02",X"2C",X"63",X"01",X"00",X"04",X"01",X"06",X"00",X"00",X"00",X"02",X"03",X"04",X"02",X"07",
		X"0A",X"04",X"02",X"0B",X"10",X"03",X"02",X"14",X"19",X"02",X"04",X"1A",X"20",X"01",X"02",X"02",
		X"02",X"01",X"01",X"02",X"02",X"35",X"27",X"01",X"02",X"2B",X"63",X"01",X"00",X"02",X"01",X"04",
		X"01",X"02",X"05",X"63",X"00",X"00",X"02",X"01",X"04",X"04",X"02",X"05",X"10",X"05",X"02",X"11",
		X"13",X"03",X"02",X"14",X"19",X"04",X"02",X"1A",X"63",X"05",X"00",X"04",X"01",X"04",X"00",X"00",
		X"01",X"00",X"02",X"05",X"10",X"01",X"02",X"11",X"20",X"01",X"02",X"21",X"27",X"01",X"02",X"28",
		X"63",X"01",X"00",X"04",X"01",X"05",X"00",X"00",X"01",X"00",X"01",X"02",X"06",X"10",X"02",X"02",
		X"11",X"1A",X"01",X"02",X"1B",X"20",X"01",X"02",X"21",X"2C",X"02",X"02",X"2D",X"63",X"03",X"00",
		X"02",X"11",X"20",X"02",X"02",X"21",X"63",X"01",X"00",X"04",X"11",X"20",X"05",X"03",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"04",X"02",X"02",X"21",X"63",X"03",
		X"00",X"02",X"0B",X"10",X"01",X"02",X"16",X"19",X"01",X"02",X"1B",X"63",X"01",X"00",X"02",X"0B",
		X"10",X"01",X"02",X"16",X"19",X"01",X"02",X"1B",X"20",X"01",X"02",X"21",X"27",X"04",X"02",X"28",
		X"63",X"03",X"00",X"04",X"11",X"12",X"28",X"14",X"0C",X"13",X"20",X"14",X"28",X"08",X"21",X"27",
		X"14",X"FF",X"0C",X"28",X"63",X"14",X"0A",X"00",X"0C",X"11",X"20",X"00",X"40",X"0C",X"21",X"30",
		X"40",X"C0",X"02",X"31",X"63",X"C0",X"00",X"02",X"01",X"10",X"DC",X"02",X"11",X"27",X"C0",X"08",
		X"28",X"40",X"C0",X"01",X"02",X"41",X"63",X"E6",X"02",X"01",X"63",X"06",X"06",X"01",X"63",X"00",
		X"00",X"00",X"E0",X"D8",X"D4",X"D0",X"C8",X"C0",X"B8",X"B0",X"A8",X"A0",X"A0",X"A0",X"A8",X"A0",
		X"9C",X"9A",X"98",X"04",X"01",X"10",X"0A",X"0C",X"0F",X"11",X"14",X"16",X"14",X"18",X"1B",X"1D",
		X"1B",X"18",X"1A",X"1C",X"1E",X"1B",X"08",X"11",X"1A",X"14",X"01",X"02",X"1B",X"27",X"1B",X"08",
		X"28",X"30",X"1D",X"01",X"08",X"31",X"40",X"1F",X"01",X"08",X"41",X"50",X"23",X"01",X"08",X"51",
		X"63",X"2B",X"01",X"02",X"01",X"14",X"02",X"02",X"15",X"20",X"02",X"02",X"21",X"63",X"03",X"02",
		X"3C",X"63",X"40",X"00",X"06",X"01",X"63",X"07",X"0B",X"19",X"24",X"53",X"0B",X"24",X"19",X"53",
		X"87",X"24",X"19",X"53",X"07",X"87",X"24",X"EF",X"95",X"6D",X"01",X"E3",X"95",X"B3",X"00",X"FA",
		X"93",X"19",X"01",X"07",X"94",X"1A",X"01",X"CD",X"94",X"29",X"01",X"D6",X"94",X"2E",X"01",X"20",
		X"95",X"2A",X"01",X"29",X"95",X"2F",X"01",X"EB",X"94",X"2B",X"01",X"03",X"95",X"30",X"01",X"89",
		X"94",X"2C",X"01",X"A5",X"94",X"31",X"01",X"41",X"95",X"2D",X"01",X"4E",X"95",X"32",X"01",X"5D",
		X"94",X"57",X"01",X"69",X"94",X"47",X"01",X"75",X"94",X"4B",X"01",X"81",X"94",X"4C",X"01",X"98",
		X"95",X"1C",X"01",X"B3",X"95",X"5B",X"01",X"9C",X"95",X"5A",X"01",X"63",X"95",X"B2",X"00",X"F4",
		X"95",X"5D",X"01",X"4D",X"94",X"63",X"01",X"49",X"94",X"20",X"01",X"1B",X"94",X"60",X"01",X"78",
		X"95",X"59",X"01",X"87",X"95",X"5F",X"01",X"AE",X"5E",X"01",X"BD",X"90",X"96",X"48",X"BD",X"8F",
		X"96",X"48",X"60",X"AE",X"5E",X"01",X"BD",X"9E",X"96",X"48",X"BD",X"9D",X"96",X"48",X"60",X"00",
		X"00",X"C3",X"96",X"B6",X"96",X"AA",X"96",X"E1",X"96",X"DA",X"96",X"FF",X"96",X"00",X"00",X"C7",
		X"96",X"CA",X"96",X"CA",X"96",X"C6",X"96",X"C7",X"96",X"C6",X"96",X"A5",X"2B",X"38",X"E9",X"01",
		X"29",X"0F",X"18",X"69",X"01",X"10",X"02",X"A5",X"2B",X"84",X"29",X"88",X"88",X"38",X"F1",X"2C",
		X"18",X"65",X"29",X"A8",X"B1",X"2C",X"60",X"C8",X"C8",X"C8",X"60",X"B1",X"2C",X"88",X"38",X"F1",
		X"2C",X"85",X"29",X"98",X"38",X"65",X"29",X"A8",X"C8",X"C8",X"60",X"B1",X"2C",X"18",X"6D",X"60",
		X"01",X"60",X"20",X"F4",X"96",X"AA",X"B1",X"2C",X"C8",X"E0",X"00",X"F0",X"06",X"18",X"71",X"2C",
		X"CA",X"D0",X"FA",X"60",X"A5",X"2B",X"84",X"29",X"88",X"88",X"38",X"F1",X"2C",X"C8",X"C8",X"60",
		X"20",X"F4",X"96",X"29",X"01",X"F0",X"01",X"C8",X"B1",X"2C",X"60",X"20",X"49",X"97",X"20",X"3F",
		X"A2",X"20",X"3A",X"A8",X"20",X"A2",X"98",X"20",X"1E",X"9B",X"20",X"8F",X"A1",X"20",X"A6",X"A2",
		X"20",X"54",X"A4",X"20",X"16",X"A4",X"4C",X"04",X"A5",X"AD",X"23",X"01",X"29",X"7F",X"8D",X"23",
		X"01",X"20",X"49",X"97",X"20",X"F8",X"97",X"20",X"16",X"A4",X"20",X"3F",X"A2",X"20",X"8F",X"A1",
		X"AD",X"01",X"02",X"10",X"03",X"20",X"04",X"A5",X"60",X"AD",X"01",X"02",X"10",X"01",X"60",X"A2",
		X"00",X"A5",X"05",X"30",X"06",X"20",X"C5",X"97",X"B8",X"50",X"15",X"A5",X"50",X"10",X"09",X"C9",
		X"E1",X"B0",X"02",X"A9",X"E1",X"B8",X"50",X"06",X"C9",X"1F",X"90",X"02",X"A9",X"1F",X"86",X"50",
		X"85",X"2B",X"49",X"FF",X"38",X"65",X"51",X"85",X"2C",X"AE",X"11",X"01",X"F0",X"1F",X"C9",X"F0",
		X"90",X"04",X"A9",X"EF",X"85",X"2C",X"45",X"2B",X"10",X"13",X"A5",X"2C",X"45",X"51",X"10",X"0D",
		X"A5",X"51",X"30",X"05",X"A9",X"00",X"B8",X"50",X"02",X"A9",X"EF",X"85",X"2C",X"A5",X"2C",X"4A",
		X"4A",X"4A",X"4A",X"85",X"2A",X"18",X"69",X"01",X"29",X"0F",X"85",X"2B",X"A5",X"2A",X"CD",X"00",
		X"02",X"F0",X"03",X"20",X"B5",X"CC",X"A5",X"2A",X"8D",X"00",X"02",X"A5",X"2B",X"8D",X"01",X"02",
		X"A5",X"2C",X"85",X"51",X"60",X"A9",X"FF",X"85",X"29",X"85",X"2A",X"AE",X"1C",X"01",X"BD",X"DF",
		X"02",X"F0",X"08",X"C5",X"29",X"B0",X"04",X"85",X"29",X"86",X"2A",X"CA",X"10",X"F0",X"A6",X"2A",
		X"30",X"15",X"BD",X"B9",X"02",X"AC",X"00",X"02",X"20",X"A6",X"A7",X"A8",X"F0",X"09",X"30",X"05",
		X"A9",X"F7",X"B8",X"50",X"02",X"A9",X"09",X"60",X"AD",X"01",X"02",X"10",X"01",X"60",X"AD",X"06",
		X"01",X"30",X"01",X"60",X"AD",X"02",X"02",X"C9",X"10",X"D0",X"03",X"20",X"EE",X"CC",X"AD",X"07",
		X"01",X"18",X"6D",X"04",X"01",X"8D",X"07",X"01",X"AD",X"02",X"02",X"6D",X"05",X"01",X"8D",X"02",
		X"02",X"B0",X"02",X"C9",X"F0",X"90",X"0C",X"A9",X"0E",X"85",X"00",X"20",X"F2",X"CC",X"A9",X"FF",
		X"8D",X"02",X"02",X"AD",X"02",X"02",X"C9",X"50",X"90",X"08",X"AD",X"15",X"01",X"D0",X"03",X"20",
		X"BD",X"A7",X"A5",X"5C",X"18",X"6D",X"04",X"01",X"85",X"5C",X"A5",X"5F",X"6D",X"05",X"01",X"90",
		X"02",X"E6",X"5B",X"C5",X"5F",X"F0",X"03",X"EE",X"14",X"01",X"85",X"5F",X"A5",X"9F",X"0A",X"0A",
		X"C9",X"30",X"90",X"02",X"A9",X"30",X"18",X"69",X"20",X"18",X"6D",X"04",X"01",X"8D",X"04",X"01",
		X"AD",X"05",X"01",X"69",X"00",X"8D",X"05",X"01",X"AD",X"02",X"02",X"C9",X"F0",X"B0",X"22",X"A2",
		X"0F",X"BD",X"AC",X"03",X"F0",X"18",X"EC",X"00",X"02",X"D0",X"13",X"CD",X"02",X"02",X"B0",X"0E",
		X"20",X"06",X"CD",X"20",X"47",X"A3",X"A9",X"00",X"8D",X"15",X"01",X"20",X"8F",X"92",X"CA",X"10",
		X"E0",X"60",X"A0",X"00",X"8C",X"4F",X"01",X"AD",X"08",X"01",X"18",X"6D",X"09",X"01",X"CD",X"1C",
		X"01",X"90",X"04",X"F0",X"02",X"A0",X"FF",X"AD",X"25",X"01",X"F0",X"02",X"A0",X"FF",X"84",X"2F",
		X"A2",X"3F",X"BD",X"43",X"02",X"F0",X"52",X"24",X"2F",X"30",X"23",X"38",X"E9",X"01",X"9D",X"43",
		X"02",X"D0",X"06",X"20",X"23",X"99",X"B8",X"50",X"15",X"C9",X"3F",X"D0",X"11",X"BC",X"03",X"02",
		X"AD",X"4F",X"01",X"0D",X"4F",X"01",X"39",X"38",X"CA",X"F0",X"03",X"FE",X"43",X"02",X"BD",X"43",
		X"02",X"C9",X"40",X"90",X"14",X"A5",X"03",X"29",X"01",X"D0",X"0B",X"BD",X"03",X"02",X"18",X"69",
		X"01",X"29",X"0F",X"9D",X"03",X"02",X"B8",X"50",X"10",X"C9",X"20",X"90",X"0C",X"BC",X"03",X"02",
		X"B9",X"38",X"CA",X"0D",X"4F",X"01",X"8D",X"4F",X"01",X"CA",X"10",X"A6",X"AD",X"4F",X"01",X"8D",
		X"50",X"01",X"60",X"A9",X"F0",X"85",X"29",X"BD",X"03",X"02",X"85",X"2A",X"86",X"35",X"20",X"A5",
		X"99",X"A6",X"35",X"A5",X"29",X"F0",X"0E",X"20",X"4D",X"99",X"F0",X"09",X"CE",X"AB",X"03",X"A9",
		X"00",X"9D",X"43",X"02",X"60",X"A9",X"FF",X"85",X"2F",X"FE",X"43",X"02",X"60",X"84",X"36",X"AC",
		X"1C",X"01",X"B9",X"DF",X"02",X"D0",X"46",X"A5",X"29",X"99",X"DF",X"02",X"A5",X"2A",X"C9",X"0F",
		X"D0",X"0A",X"2C",X"11",X"01",X"10",X"05",X"AD",X"CA",X"60",X"29",X"0E",X"99",X"B9",X"02",X"18",
		X"69",X"01",X"29",X"0F",X"99",X"CC",X"02",X"A9",X"00",X"99",X"A6",X"02",X"A5",X"2C",X"99",X"8A",
		X"02",X"A5",X"2D",X"99",X"91",X"02",X"EE",X"08",X"01",X"A5",X"2B",X"99",X"83",X"02",X"A4",X"36",
		X"29",X"07",X"86",X"36",X"AA",X"FE",X"42",X"01",X"A6",X"36",X"A9",X"10",X"60",X"88",X"10",X"B2",
		X"A4",X"36",X"A9",X"00",X"60",X"A9",X"00",X"A2",X"04",X"9D",X"3D",X"01",X"CA",X"10",X"FA",X"A2",
		X"04",X"BD",X"2E",X"01",X"38",X"FD",X"42",X"01",X"90",X"03",X"9D",X"3D",X"01",X"CA",X"10",X"F1",
		X"AC",X"1C",X"01",X"B9",X"DF",X"02",X"F0",X"14",X"B9",X"8A",X"02",X"29",X"03",X"F0",X"0D",X"AA",
		X"E0",X"03",X"D0",X"02",X"A2",X"05",X"DE",X"3C",X"01",X"DE",X"3C",X"01",X"88",X"10",X"E4",X"A2",
		X"04",X"AD",X"1C",X"01",X"18",X"69",X"01",X"38",X"FD",X"42",X"01",X"CA",X"10",X"F9",X"A2",X"04",
		X"DD",X"3D",X"01",X"B0",X"03",X"9D",X"3D",X"01",X"CA",X"10",X"F5",X"A2",X"04",X"A0",X"00",X"BD",
		X"3D",X"01",X"F0",X"01",X"C8",X"CA",X"10",X"F7",X"98",X"F0",X"77",X"88",X"D0",X"18",X"A2",X"04",
		X"BD",X"3D",X"01",X"F0",X"0B",X"BD",X"29",X"01",X"F0",X"06",X"20",X"87",X"9A",X"F0",X"01",X"60",
		X"CA",X"10",X"ED",X"B8",X"50",X"5C",X"84",X"61",X"A2",X"04",X"BD",X"3D",X"01",X"F0",X"0E",X"BD",
		X"42",X"01",X"DD",X"29",X"01",X"B0",X"06",X"20",X"87",X"9A",X"F0",X"01",X"60",X"CA",X"10",X"EA",
		X"AD",X"40",X"01",X"F0",X"1C",X"AD",X"3F",X"01",X"F0",X"17",X"A4",X"2A",X"B9",X"AC",X"03",X"D0",
		X"02",X"A9",X"FF",X"A2",X"03",X"C9",X"CC",X"B0",X"02",X"A2",X"02",X"20",X"87",X"9A",X"F0",X"01",
		X"60",X"AD",X"DA",X"60",X"29",X"03",X"AA",X"E8",X"A0",X"04",X"BD",X"29",X"01",X"F0",X"0B",X"BD",
		X"3D",X"01",X"F0",X"06",X"20",X"87",X"9A",X"F0",X"01",X"60",X"CA",X"10",X"02",X"A2",X"04",X"88",
		X"10",X"E8",X"A9",X"00",X"85",X"29",X"60",X"8A",X"0A",X"A8",X"B9",X"94",X"9A",X"48",X"B9",X"93",
		X"9A",X"48",X"60",X"9C",X"9A",X"A8",X"9A",X"BA",X"9A",X"B6",X"9A",X"B2",X"9A",X"AD",X"02",X"9B",
		X"85",X"2C",X"AD",X"5D",X"01",X"A0",X"00",X"F0",X"4D",X"AD",X"03",X"9B",X"0D",X"6D",X"01",X"A0",
		X"01",X"D0",X"3E",X"A0",X"04",X"D0",X"37",X"A0",X"03",X"D0",X"33",X"AD",X"CA",X"60",X"29",X"03",
		X"A8",X"A9",X"04",X"85",X"2B",X"86",X"39",X"C6",X"2B",X"10",X"05",X"A6",X"39",X"A9",X"00",X"60",
		X"88",X"10",X"02",X"A0",X"03",X"BE",X"49",X"01",X"E0",X"03",X"D0",X"02",X"A2",X"05",X"BD",X"3C",
		X"01",X"F0",X"E4",X"A6",X"39",X"B9",X"49",X"01",X"09",X"40",X"A0",X"02",X"D0",X"03",X"B9",X"02",
		X"9B",X"85",X"2C",X"B9",X"FD",X"9A",X"84",X"2B",X"85",X"2D",X"A5",X"29",X"60",X"07",X"72",X"07",
		X"00",X"61",X"40",X"00",X"41",X"40",X"00",X"84",X"36",X"A5",X"29",X"C9",X"20",X"A5",X"2B",X"B0",
		X"07",X"A8",X"20",X"EE",X"9A",X"B8",X"50",X"03",X"20",X"88",X"9A",X"A4",X"36",X"60",X"AD",X"01",
		X"02",X"30",X"33",X"AE",X"1C",X"01",X"86",X"37",X"A6",X"37",X"BD",X"DF",X"02",X"F0",X"23",X"A9",
		X"01",X"8D",X"0A",X"01",X"BD",X"91",X"02",X"8D",X"0B",X"01",X"AD",X"0B",X"01",X"A8",X"B9",X"F7",
		X"A0",X"20",X"98",X"9B",X"EE",X"0B",X"01",X"AD",X"0A",X"01",X"D0",X"EE",X"AD",X"0B",X"01",X"9D",
		X"91",X"02",X"C6",X"37",X"10",X"D2",X"AD",X"48",X"01",X"18",X"6D",X"47",X"01",X"A8",X"4D",X"48",
		X"01",X"8C",X"48",X"01",X"10",X"16",X"98",X"10",X"06",X"20",X"06",X"CD",X"B8",X"50",X"0D",X"AD",
		X"43",X"01",X"F0",X"08",X"AD",X"01",X"02",X"30",X"03",X"20",X"02",X"CD",X"AD",X"48",X"01",X"30",
		X"07",X"C9",X"0F",X"B0",X"07",X"B8",X"50",X"0F",X"C9",X"C1",X"B0",X"0B",X"AD",X"47",X"01",X"49",
		X"FF",X"18",X"69",X"01",X"8D",X"47",X"01",X"60",X"A8",X"B9",X"A3",X"9B",X"48",X"B9",X"A2",X"9B",
		X"48",X"60",X"C9",X"9B",X"CF",X"9B",X"ED",X"9B",X"16",X"9C",X"0B",X"9C",X"CE",X"9B",X"57",X"9C",
		X"C3",X"9F",X"DC",X"9B",X"5B",X"9E",X"81",X"9D",X"4E",X"9C",X"2E",X"9E",X"F9",X"9B",X"20",X"9C",
		X"F0",X"9E",X"47",X"9E",X"B5",X"9C",X"66",X"9D",X"3A",X"9C",X"A9",X"00",X"8D",X"0A",X"01",X"60",
		X"EE",X"0B",X"01",X"AC",X"0B",X"01",X"B9",X"F7",X"A0",X"9D",X"98",X"02",X"60",X"EE",X"0B",X"01",
		X"AC",X"0B",X"01",X"B9",X"F7",X"A0",X"A8",X"B9",X"00",X"00",X"9D",X"98",X"02",X"60",X"AD",X"0C",
		X"01",X"D0",X"06",X"EE",X"0B",X"01",X"EE",X"0B",X"01",X"60",X"EE",X"0B",X"01",X"AD",X"0C",X"01",
		X"D0",X"09",X"AC",X"0B",X"01",X"B9",X"F7",X"A0",X"8D",X"0B",X"01",X"60",X"DE",X"98",X"02",X"D0",
		X"06",X"EE",X"0B",X"01",X"B8",X"50",X"09",X"AC",X"0B",X"01",X"B9",X"F8",X"A0",X"8D",X"0B",X"01",
		X"60",X"BC",X"B9",X"02",X"B9",X"AC",X"03",X"D0",X"02",X"A9",X"FF",X"DD",X"DF",X"02",X"B0",X"05",
		X"A9",X"00",X"B8",X"50",X"02",X"A9",X"01",X"8D",X"0C",X"01",X"60",X"AD",X"47",X"01",X"0A",X"0A",
		X"18",X"6D",X"48",X"01",X"2D",X"48",X"01",X"29",X"80",X"49",X"80",X"8D",X"0C",X"01",X"60",X"BD",
		X"83",X"02",X"49",X"40",X"9D",X"83",X"02",X"60",X"BD",X"83",X"02",X"29",X"07",X"A8",X"BD",X"8A",
		X"02",X"30",X"36",X"BD",X"9F",X"02",X"18",X"79",X"60",X"01",X"9D",X"9F",X"02",X"BD",X"DF",X"02",
		X"79",X"65",X"01",X"9D",X"DF",X"02",X"CD",X"02",X"02",X"F0",X"02",X"B0",X"06",X"20",X"06",X"9D",
		X"B8",X"50",X"13",X"C9",X"20",X"B0",X"0F",X"BD",X"8A",X"02",X"29",X"03",X"F0",X"08",X"8A",X"48",
		X"A8",X"20",X"6F",X"A0",X"68",X"AA",X"B8",X"50",X"1C",X"BD",X"9F",X"02",X"38",X"F9",X"60",X"01",
		X"9D",X"9F",X"02",X"BD",X"DF",X"02",X"F9",X"65",X"01",X"9D",X"DF",X"02",X"C9",X"F0",X"90",X"05",
		X"A9",X"F2",X"9D",X"DF",X"02",X"60",X"A0",X"01",X"BD",X"8A",X"02",X"30",X"10",X"BD",X"DF",X"02",
		X"CD",X"57",X"01",X"90",X"02",X"A0",X"00",X"20",X"63",X"9C",X"B8",X"50",X"17",X"20",X"99",X"9C",
		X"AC",X"AB",X"03",X"D0",X"02",X"A9",X"FF",X"CD",X"57",X"01",X"90",X"08",X"BD",X"8A",X"02",X"49",
		X"80",X"9D",X"8A",X"02",X"AD",X"48",X"01",X"30",X"1B",X"BD",X"DF",X"02",X"CD",X"57",X"01",X"B0",
		X"13",X"AD",X"00",X"02",X"DD",X"B9",X"02",X"D0",X"0B",X"AD",X"01",X"02",X"DD",X"CC",X"02",X"D0",
		X"03",X"20",X"47",X"A3",X"60",X"16",X"AD",X"02",X"02",X"9D",X"DF",X"02",X"BD",X"83",X"02",X"29",
		X"07",X"C9",X"01",X"D0",X"0E",X"AD",X"AB",X"03",X"F0",X"09",X"BD",X"8A",X"02",X"49",X"80",X"9D",
		X"8A",X"02",X"60",X"BD",X"83",X"02",X"10",X"04",X"FE",X"DF",X"02",X"60",X"CE",X"08",X"01",X"AD",
		X"09",X"01",X"C9",X"01",X"F0",X"06",X"20",X"67",X"9D",X"B8",X"50",X"22",X"A0",X"06",X"B9",X"DF",
		X"02",X"F0",X"0E",X"84",X"38",X"E4",X"38",X"F0",X"08",X"B9",X"DF",X"02",X"CD",X"02",X"02",X"F0",
		X"03",X"88",X"10",X"EA",X"B9",X"83",X"02",X"29",X"40",X"49",X"40",X"9D",X"83",X"02",X"A9",X"41",
		X"8D",X"0B",X"01",X"EE",X"09",X"01",X"60",X"BD",X"B9",X"02",X"A8",X"AD",X"00",X"02",X"20",X"A6",
		X"A7",X"0A",X"BD",X"83",X"02",X"B0",X"05",X"09",X"40",X"B8",X"50",X"02",X"29",X"BF",X"9D",X"83",
		X"02",X"60",X"BC",X"CC",X"02",X"BD",X"83",X"02",X"29",X"40",X"D0",X"04",X"C8",X"B8",X"50",X"01",
		X"88",X"98",X"29",X"0F",X"09",X"80",X"9D",X"CC",X"02",X"BD",X"83",X"02",X"29",X"07",X"C9",X"04",
		X"D0",X"4C",X"BD",X"CC",X"02",X"29",X"07",X"D0",X"42",X"BD",X"CC",X"02",X"29",X"08",X"F0",X"0B",
		X"BD",X"B9",X"02",X"18",X"69",X"01",X"29",X"0F",X"9D",X"B9",X"02",X"BD",X"83",X"02",X"29",X"7F",
		X"9D",X"83",X"02",X"A9",X"20",X"9D",X"CC",X"02",X"BD",X"8A",X"02",X"49",X"80",X"9D",X"8A",X"02",
		X"AD",X"AB",X"03",X"D0",X"16",X"BD",X"DF",X"02",X"CD",X"02",X"02",X"D0",X"06",X"20",X"81",X"9F",
		X"B8",X"50",X"08",X"BD",X"8A",X"02",X"29",X"80",X"9D",X"8A",X"02",X"B8",X"50",X"38",X"BC",X"B9",
		X"02",X"BD",X"83",X"02",X"49",X"40",X"20",X"D7",X"9E",X"DD",X"CC",X"02",X"D0",X"28",X"BD",X"83",
		X"02",X"29",X"7F",X"9D",X"83",X"02",X"29",X"40",X"D0",X"11",X"BD",X"B9",X"02",X"9D",X"CC",X"02",
		X"38",X"E9",X"01",X"29",X"0F",X"9D",X"B9",X"02",X"B8",X"50",X"0B",X"BD",X"B9",X"02",X"18",X"69",
		X"01",X"29",X"0F",X"9D",X"CC",X"02",X"BD",X"83",X"02",X"29",X"80",X"8D",X"0C",X"01",X"60",X"BD",
		X"83",X"02",X"30",X"13",X"BD",X"B9",X"02",X"CD",X"00",X"02",X"D0",X"0B",X"BD",X"CC",X"02",X"CD",
		X"01",X"02",X"D0",X"03",X"20",X"3A",X"A3",X"60",X"BD",X"DF",X"02",X"CD",X"02",X"02",X"D0",X"0B",
		X"BD",X"B9",X"02",X"CD",X"00",X"02",X"D0",X"03",X"20",X"43",X"A3",X"60",X"20",X"AB",X"9E",X"BD",
		X"83",X"02",X"09",X"80",X"9D",X"83",X"02",X"29",X"07",X"C9",X"04",X"D0",X"1F",X"BD",X"83",X"02",
		X"29",X"40",X"D0",X"05",X"A9",X"81",X"B8",X"50",X"0D",X"BD",X"B9",X"02",X"38",X"E9",X"01",X"29",
		X"0F",X"9D",X"B9",X"02",X"A9",X"87",X"9D",X"CC",X"02",X"B8",X"50",X"1E",X"BD",X"83",X"02",X"29",
		X"40",X"F0",X"0B",X"BD",X"B9",X"02",X"18",X"69",X"01",X"29",X"0F",X"9D",X"B9",X"02",X"BD",X"83",
		X"02",X"BC",X"B9",X"02",X"20",X"D7",X"9E",X"9D",X"CC",X"02",X"60",X"AD",X"11",X"01",X"F0",X"26",
		X"BD",X"83",X"02",X"29",X"40",X"F0",X"12",X"BD",X"B9",X"02",X"C9",X"0E",X"90",X"08",X"BD",X"83",
		X"02",X"29",X"BF",X"9D",X"83",X"02",X"B8",X"50",X"0D",X"BD",X"B9",X"02",X"D0",X"08",X"BD",X"83",
		X"02",X"09",X"40",X"9D",X"83",X"02",X"60",X"29",X"40",X"F0",X"10",X"88",X"98",X"29",X"0F",X"A8",
		X"B9",X"EE",X"03",X"18",X"69",X"08",X"29",X"0F",X"B8",X"50",X"03",X"B9",X"EE",X"03",X"09",X"80",
		X"60",X"A0",X"04",X"BD",X"8A",X"02",X"30",X"4B",X"BD",X"9F",X"02",X"18",X"6D",X"64",X"01",X"9D",
		X"9F",X"02",X"BD",X"DF",X"02",X"6D",X"69",X"01",X"9D",X"DF",X"02",X"CD",X"02",X"02",X"B0",X"09",
		X"AD",X"02",X"02",X"9D",X"DF",X"02",X"B8",X"50",X"11",X"AC",X"AB",X"03",X"F0",X"0B",X"A4",X"9F",
		X"C0",X"11",X"B0",X"02",X"C9",X"20",X"B8",X"50",X"01",X"60",X"B0",X"11",X"AD",X"59",X"01",X"10",
		X"06",X"20",X"81",X"9F",X"B8",X"50",X"03",X"20",X"8A",X"9F",X"B8",X"50",X"03",X"20",X"5F",X"9F",
		X"B8",X"50",X"1B",X"20",X"99",X"9C",X"C9",X"80",X"90",X"11",X"2C",X"59",X"01",X"50",X"06",X"20",
		X"81",X"9F",X"B8",X"50",X"03",X"20",X"8A",X"9F",X"B8",X"50",X"03",X"20",X"5F",X"9F",X"60",X"BD",
		X"DF",X"02",X"29",X"20",X"F0",X"1A",X"AD",X"DA",X"60",X"CD",X"5F",X"01",X"90",X"12",X"2C",X"59",
		X"01",X"50",X"0A",X"8A",X"4A",X"90",X"13",X"20",X"81",X"9F",X"B8",X"50",X"03",X"20",X"8A",X"9F",
		X"60",X"20",X"67",X"9D",X"20",X"4F",X"9C",X"4C",X"99",X"9F",X"BD",X"83",X"02",X"29",X"BF",X"2C",
		X"CA",X"60",X"50",X"02",X"09",X"40",X"9D",X"83",X"02",X"AD",X"11",X"01",X"F0",X"1E",X"BD",X"83",
		X"02",X"29",X"40",X"D0",X"0A",X"BD",X"B9",X"02",X"C9",X"0F",X"B0",X"08",X"B8",X"50",X"0D",X"BD",
		X"B9",X"02",X"D0",X"08",X"BD",X"83",X"02",X"49",X"40",X"9D",X"83",X"02",X"A9",X"66",X"8D",X"0B",
		X"01",X"4C",X"5F",X"9E",X"A9",X"01",X"8D",X"0C",X"01",X"BC",X"B9",X"02",X"B9",X"AC",X"03",X"D0",
		X"05",X"A9",X"F1",X"99",X"AC",X"03",X"BD",X"DF",X"02",X"D9",X"AC",X"03",X"B0",X"08",X"99",X"AC",
		X"03",X"A9",X"80",X"99",X"9A",X"03",X"BD",X"DF",X"02",X"C9",X"20",X"B0",X"10",X"BD",X"8A",X"02",
		X"09",X"80",X"9D",X"8A",X"02",X"A9",X"20",X"9D",X"DF",X"02",X"B8",X"50",X"2A",X"C9",X"F2",X"90",
		X"26",X"20",X"28",X"A0",X"A9",X"F0",X"9D",X"DF",X"02",X"AD",X"AB",X"03",X"D0",X"19",X"BD",X"8A",
		X"02",X"29",X"FC",X"09",X"01",X"9D",X"8A",X"02",X"BD",X"83",X"02",X"29",X"F8",X"09",X"02",X"9D",
		X"83",X"02",X"A9",X"00",X"8D",X"0C",X"01",X"60",X"A9",X"00",X"85",X"2D",X"A9",X"0F",X"8D",X"40",
		X"01",X"AD",X"DA",X"60",X"29",X"0F",X"A8",X"C0",X"0F",X"D0",X"05",X"AD",X"11",X"01",X"D0",X"0F",
		X"B9",X"AC",X"03",X"D0",X"02",X"A9",X"FF",X"C5",X"2D",X"90",X"04",X"85",X"2D",X"84",X"29",X"88",
		X"10",X"02",X"A0",X"0F",X"CE",X"40",X"01",X"10",X"DE",X"A5",X"29",X"9D",X"B9",X"02",X"18",X"69",
		X"01",X"29",X"0F",X"9D",X"CC",X"02",X"BD",X"8A",X"02",X"29",X"7F",X"9D",X"8A",X"02",X"60",X"B9",
		X"DF",X"02",X"85",X"29",X"CD",X"02",X"02",X"D0",X"0F",X"B9",X"83",X"02",X"29",X"07",X"C9",X"04",
		X"F0",X"06",X"CE",X"09",X"01",X"B8",X"50",X"03",X"CE",X"08",X"01",X"A9",X"00",X"99",X"DF",X"02",
		X"B9",X"83",X"02",X"29",X"07",X"86",X"35",X"AA",X"DE",X"42",X"01",X"A6",X"35",X"B9",X"8A",X"02",
		X"29",X"03",X"F0",X"52",X"38",X"E9",X"01",X"C9",X"02",X"D0",X"02",X"A9",X"04",X"85",X"2B",X"B9",
		X"B9",X"02",X"38",X"E9",X"01",X"29",X"0F",X"C9",X"0F",X"90",X"07",X"2C",X"11",X"01",X"10",X"02",
		X"A9",X"00",X"85",X"2A",X"20",X"07",X"9B",X"A5",X"2D",X"8D",X"0B",X"01",X"CE",X"0B",X"01",X"A9",
		X"00",X"8D",X"0A",X"01",X"20",X"4D",X"99",X"F0",X"1D",X"A5",X"2A",X"18",X"69",X"02",X"29",X"0F",
		X"C9",X"0F",X"D0",X"07",X"2C",X"11",X"01",X"10",X"02",X"A9",X"0E",X"85",X"2A",X"A5",X"2B",X"09",
		X"40",X"85",X"2B",X"20",X"4D",X"99",X"60",X"0C",X"0E",X"1A",X"06",X"00",X"06",X"FF",X"0C",X"00",
		X"06",X"06",X"02",X"08",X"0C",X"00",X"08",X"0C",X"12",X"00",X"14",X"04",X"06",X"11",X"06",X"0A",
		X"0C",X"00",X"12",X"00",X"14",X"0C",X"04",X"06",X"1B",X"06",X"18",X"0C",X"00",X"02",X"02",X"12",
		X"00",X"14",X"0C",X"04",X"06",X"28",X"00",X"08",X"27",X"16",X"02",X"03",X"12",X"00",X"14",X"0C",
		X"04",X"06",X"35",X"00",X"08",X"34",X"16",X"06",X"23",X"02",X"04",X"18",X"00",X"08",X"43",X"12",
		X"00",X"10",X"B3",X"14",X"1A",X"41",X"08",X"4B",X"06",X"48",X"00",X"0C",X"1C",X"1A",X"52",X"12",
		X"00",X"0C",X"14",X"1A",X"52",X"00",X"06",X"5A",X"1E",X"20",X"00",X"06",X"60",X"00",X"02",X"03",
		X"20",X"00",X"08",X"68",X"14",X"1A",X"60",X"06",X"65",X"10",X"B2",X"22",X"00",X"08",X"73",X"26",
		X"1A",X"7E",X"22",X"00",X"06",X"77",X"24",X"12",X"00",X"14",X"1A",X"71",X"06",X"80",X"24",X"16",
		X"12",X"00",X"0C",X"14",X"04",X"06",X"89",X"02",X"04",X"00",X"0C",X"08",X"91",X"06",X"86",X"A2",
		X"0B",X"86",X"37",X"A6",X"37",X"BD",X"D3",X"02",X"F0",X"45",X"E0",X"08",X"B0",X"22",X"69",X"09",
		X"BC",X"F2",X"02",X"F0",X"03",X"38",X"E9",X"04",X"9D",X"D3",X"02",X"20",X"FA",X"A1",X"BD",X"D3",
		X"02",X"C9",X"F0",X"90",X"08",X"CE",X"35",X"01",X"A9",X"00",X"9D",X"D3",X"02",X"B8",X"50",X"1F",
		X"BD",X"E6",X"02",X"18",X"6D",X"20",X"01",X"9D",X"E6",X"02",X"BD",X"D3",X"02",X"6D",X"18",X"01",
		X"CD",X"02",X"02",X"B0",X"07",X"C6",X"A6",X"20",X"E4",X"A1",X"A9",X"00",X"9D",X"D3",X"02",X"C6",
		X"37",X"10",X"B0",X"60",X"AD",X"00",X"02",X"DD",X"AD",X"02",X"D0",X"0D",X"AD",X"01",X"02",X"30",
		X"08",X"20",X"4B",X"A3",X"A9",X"81",X"8D",X"01",X"02",X"60",X"BC",X"AD",X"02",X"B9",X"AC",X"03",
		X"F0",X"3C",X"BD",X"D3",X"02",X"D9",X"AC",X"03",X"90",X"25",X"C9",X"F0",X"90",X"02",X"A9",X"00",
		X"99",X"AC",X"03",X"FE",X"F2",X"02",X"A9",X"C0",X"99",X"9A",X"03",X"20",X"F6",X"CC",X"A2",X"FF",
		X"A9",X"00",X"85",X"2A",X"85",X"2B",X"A9",X"01",X"85",X"29",X"20",X"6C",X"CA",X"A6",X"37",X"BD",
		X"F2",X"02",X"C9",X"02",X"90",X"08",X"A9",X"00",X"9D",X"D3",X"02",X"CE",X"35",X"01",X"60",X"AD",
		X"01",X"02",X"30",X"61",X"A5",X"05",X"30",X"28",X"AD",X"06",X"01",X"85",X"29",X"A2",X"0A",X"BD",
		X"DB",X"02",X"F0",X"14",X"BD",X"B5",X"02",X"38",X"ED",X"00",X"02",X"10",X"05",X"49",X"FF",X"18",
		X"69",X"01",X"C9",X"02",X"B0",X"02",X"E6",X"29",X"CA",X"10",X"E4",X"A5",X"29",X"B8",X"50",X"04",
		X"A5",X"4D",X"29",X"10",X"F0",X"2F",X"A2",X"07",X"BD",X"D3",X"02",X"D0",X"25",X"EE",X"35",X"01",
		X"AD",X"02",X"02",X"9D",X"D3",X"02",X"AD",X"00",X"02",X"9D",X"AD",X"02",X"AD",X"01",X"02",X"9D",
		X"C0",X"02",X"A9",X"00",X"9D",X"F2",X"02",X"20",X"EA",X"CC",X"AD",X"02",X"02",X"20",X"63",X"A4",
		X"A2",X"00",X"CA",X"10",X"D3",X"60",X"AD",X"01",X"02",X"30",X"58",X"A2",X"06",X"BD",X"DF",X"02",
		X"F0",X"4E",X"C9",X"30",X"90",X"4A",X"BD",X"8A",X"02",X"29",X"40",X"F0",X"43",X"DE",X"A6",X"02",
		X"10",X"3E",X"FE",X"A6",X"02",X"BD",X"83",X"02",X"29",X"80",X"D0",X"34",X"AD",X"CA",X"60",X"A4",
		X"A6",X"D9",X"04",X"A3",X"90",X"2A",X"AC",X"1A",X"01",X"B9",X"DB",X"02",X"D0",X"1F",X"BD",X"DF",
		X"02",X"99",X"DB",X"02",X"BD",X"B9",X"02",X"99",X"B5",X"02",X"BD",X"CC",X"02",X"99",X"C8",X"02",
		X"AD",X"19",X"01",X"9D",X"A6",X"02",X"20",X"BD",X"CC",X"E6",X"A6",X"A0",X"00",X"88",X"10",X"D9",
		X"CA",X"10",X"AA",X"60",X"00",X"E0",X"F0",X"FA",X"FF",X"86",X"37",X"A9",X"FF",X"9D",X"F2",X"02",
		X"98",X"38",X"E9",X"04",X"A8",X"B9",X"B9",X"02",X"85",X"2D",X"AD",X"DA",X"60",X"29",X"07",X"C9",
		X"03",X"90",X"02",X"A9",X"00",X"48",X"18",X"69",X"02",X"20",X"CA",X"A3",X"20",X"6F",X"A0",X"68",
		X"18",X"69",X"05",X"AA",X"20",X"6C",X"CA",X"A6",X"37",X"60",X"A9",X"05",X"20",X"52",X"A3",X"CE",
		X"01",X"02",X"60",X"A9",X"09",X"D0",X"06",X"A9",X"07",X"D0",X"02",X"A9",X"FF",X"8D",X"3B",X"01",
		X"A9",X"01",X"85",X"2C",X"AD",X"02",X"02",X"85",X"29",X"AD",X"00",X"02",X"85",X"2D",X"20",X"B0",
		X"CC",X"20",X"D6",X"A3",X"A9",X"81",X"8D",X"01",X"02",X"A9",X"01",X"8D",X"3C",X"01",X"60",X"20",
		X"C1",X"CC",X"B9",X"DB",X"02",X"85",X"29",X"B9",X"B5",X"02",X"85",X"2D",X"A9",X"00",X"20",X"D4",
		X"A3",X"A9",X"00",X"99",X"DB",X"02",X"C6",X"A6",X"A9",X"FF",X"9D",X"F2",X"02",X"60",X"A9",X"FF",
		X"9D",X"F2",X"02",X"98",X"38",X"E9",X"04",X"A8",X"B9",X"83",X"02",X"29",X"C0",X"C9",X"C0",X"F0",
		X"06",X"B9",X"B9",X"02",X"B8",X"50",X"08",X"B9",X"B9",X"02",X"38",X"E9",X"01",X"29",X"0F",X"85",
		X"2D",X"A9",X"00",X"20",X"CA",X"A3",X"20",X"6F",X"A0",X"B9",X"83",X"02",X"29",X"07",X"A8",X"BE",
		X"C5",X"A3",X"4C",X"6C",X"CA",X"01",X"02",X"03",X"04",X"01",X"48",X"20",X"C1",X"CC",X"B9",X"DF",
		X"02",X"85",X"29",X"68",X"85",X"2C",X"86",X"35",X"84",X"36",X"A9",X"00",X"85",X"2A",X"85",X"2B",
		X"A2",X"07",X"BD",X"0A",X"03",X"F0",X"13",X"BD",X"12",X"03",X"C5",X"2A",X"90",X"04",X"85",X"2A",
		X"86",X"2B",X"CA",X"10",X"ED",X"CE",X"16",X"01",X"A6",X"2B",X"A9",X"00",X"9D",X"12",X"03",X"A5",
		X"2C",X"9D",X"02",X"03",X"A5",X"29",X"9D",X"0A",X"03",X"A5",X"2D",X"9D",X"FA",X"02",X"EE",X"16",
		X"01",X"A6",X"35",X"A4",X"36",X"60",X"AD",X"16",X"01",X"F0",X"2C",X"A9",X"00",X"8D",X"16",X"01",
		X"A2",X"07",X"BD",X"0A",X"03",X"F0",X"1D",X"BD",X"12",X"03",X"BC",X"02",X"03",X"18",X"79",X"4E",
		X"A4",X"9D",X"12",X"03",X"D9",X"48",X"A4",X"90",X"08",X"A9",X"00",X"9D",X"0A",X"03",X"B8",X"50",
		X"03",X"EE",X"16",X"01",X"CA",X"10",X"DB",X"60",X"10",X"15",X"20",X"20",X"20",X"10",X"03",X"01",
		X"03",X"03",X"03",X"03",X"A2",X"07",X"BD",X"D3",X"02",X"F0",X"03",X"20",X"63",X"A4",X"CA",X"10",
		X"F5",X"60",X"AB",X"85",X"2E",X"A0",X"0A",X"B9",X"DB",X"02",X"F0",X"7F",X"C5",X"2E",X"90",X"05",
		X"E5",X"2E",X"B8",X"50",X"06",X"A5",X"2E",X"38",X"F9",X"DB",X"02",X"C0",X"04",X"B0",X"12",X"C5",
		X"A7",X"B0",X"0B",X"B9",X"B5",X"02",X"5D",X"AD",X"02",X"D0",X"03",X"20",X"6F",X"A3",X"B8",X"50",
		X"5A",X"48",X"84",X"38",X"B9",X"7F",X"02",X"29",X"07",X"A8",X"68",X"D9",X"51",X"01",X"B0",X"49",
		X"C0",X"04",X"D0",X"1D",X"A4",X"38",X"B9",X"DB",X"02",X"CD",X"02",X"02",X"F0",X"10",X"BD",X"AD",
		X"02",X"D9",X"B5",X"02",X"D0",X"08",X"B9",X"C8",X"02",X"10",X"03",X"20",X"09",X"A3",X"B8",X"50",
		X"28",X"A4",X"38",X"B9",X"C8",X"02",X"10",X"0A",X"B9",X"B5",X"02",X"DD",X"C0",X"02",X"F0",X"12",
		X"D0",X"08",X"B9",X"DB",X"02",X"CD",X"02",X"02",X"F0",X"0F",X"B9",X"B5",X"02",X"DD",X"AD",X"02",
		X"D0",X"07",X"86",X"37",X"20",X"8E",X"A3",X"A6",X"37",X"A4",X"38",X"88",X"30",X"03",X"4C",X"67",
		X"A4",X"BD",X"F2",X"02",X"C9",X"FF",X"D0",X"0B",X"A9",X"00",X"9D",X"D3",X"02",X"CE",X"35",X"01",
		X"9D",X"F2",X"02",X"60",X"AD",X"01",X"02",X"10",X"78",X"AD",X"35",X"01",X"05",X"A6",X"0D",X"16",
		X"01",X"D0",X"6B",X"AE",X"1C",X"01",X"BD",X"DF",X"02",X"F0",X"0E",X"18",X"69",X"0F",X"B0",X"02",
		X"C9",X"F0",X"90",X"02",X"A9",X"00",X"9D",X"DF",X"02",X"CA",X"10",X"EA",X"A6",X"3D",X"B5",X"48",
		X"C9",X"01",X"D0",X"20",X"A9",X"00",X"8D",X"0F",X"01",X"A9",X"01",X"8D",X"14",X"01",X"A5",X"5F",
		X"38",X"E9",X"20",X"85",X"5F",X"A5",X"5B",X"E9",X"00",X"85",X"5B",X"C9",X"FA",X"18",X"D0",X"01",
		X"38",X"B8",X"50",X"0D",X"AD",X"02",X"02",X"18",X"69",X"0F",X"8D",X"02",X"02",X"B0",X"02",X"C9",
		X"F0",X"90",X"1B",X"A9",X"06",X"85",X"00",X"20",X"8F",X"92",X"AD",X"08",X"01",X"18",X"6D",X"09",
		X"01",X"18",X"6D",X"AB",X"03",X"C9",X"3F",X"90",X"02",X"A9",X"3F",X"8D",X"AB",X"03",X"B8",X"50",
		X"49",X"AD",X"55",X"04",X"0D",X"1B",X"01",X"F0",X"0A",X"A9",X"17",X"C5",X"42",X"B0",X"04",X"A6",
		X"40",X"F6",X"00",X"AD",X"06",X"01",X"D0",X"32",X"AD",X"AB",X"03",X"0D",X"16",X"01",X"D0",X"15",
		X"AC",X"1C",X"01",X"B9",X"DF",X"02",X"F0",X"04",X"C9",X"11",X"B0",X"09",X"88",X"10",X"F4",X"20",
		X"CB",X"A5",X"20",X"8F",X"92",X"A5",X"4D",X"29",X"60",X"F0",X"0F",X"24",X"05",X"10",X"0B",X"A5",
		X"09",X"29",X"43",X"C9",X"40",X"D0",X"03",X"20",X"CB",X"A5",X"60",X"A9",X"20",X"85",X"00",X"AD",
		X"06",X"01",X"09",X"80",X"8D",X"06",X"01",X"A9",X"00",X"8D",X"04",X"01",X"8D",X"07",X"01",X"85",
		X"5C",X"8D",X"23",X"01",X"A9",X"02",X"8D",X"05",X"01",X"A2",X"0F",X"BD",X"AC",X"03",X"F0",X"03",
		X"EE",X"23",X"01",X"CA",X"10",X"F5",X"AD",X"23",X"01",X"F0",X"17",X"A5",X"9F",X"C9",X"07",X"B0",
		X"11",X"A9",X"1E",X"85",X"04",X"A9",X"0A",X"85",X"00",X"A9",X"20",X"85",X"02",X"A9",X"80",X"8D",
		X"23",X"01",X"A9",X"FF",X"8D",X"25",X"01",X"60",X"AD",X"0E",X"01",X"8D",X"0D",X"01",X"A2",X"0F",
		X"86",X"37",X"A6",X"37",X"BD",X"83",X"02",X"D0",X"0B",X"AD",X"0E",X"01",X"F0",X"03",X"20",X"5B",
		X"A6",X"B8",X"50",X"0B",X"20",X"A9",X"A6",X"20",X"21",X"A7",X"A9",X"FF",X"8D",X"0D",X"01",X"C6",
		X"37",X"10",X"DF",X"A5",X"03",X"29",X"01",X"D0",X"08",X"AD",X"0E",X"01",X"F0",X"03",X"CE",X"0E",
		X"01",X"AD",X"0D",X"01",X"D0",X"04",X"A9",X"12",X"85",X"00",X"60",X"A5",X"03",X"29",X"00",X"D0",
		X"39",X"A9",X"80",X"9D",X"63",X"02",X"9D",X"83",X"02",X"9D",X"A3",X"02",X"AD",X"DA",X"60",X"9D",
		X"C3",X"02",X"20",X"9B",X"A6",X"9D",X"23",X"03",X"AD",X"CA",X"60",X"9D",X"E3",X"02",X"20",X"9B",
		X"A6",X"30",X"05",X"49",X"FF",X"18",X"69",X"01",X"9D",X"43",X"03",X"AD",X"CA",X"60",X"9D",X"03",
		X"03",X"20",X"9B",X"A6",X"9D",X"63",X"03",X"20",X"C1",X"CC",X"60",X"4A",X"AD",X"DA",X"60",X"29",
		X"07",X"90",X"05",X"49",X"FF",X"18",X"69",X"01",X"60",X"BD",X"E3",X"02",X"18",X"7D",X"23",X"02",
		X"9D",X"23",X"02",X"BD",X"43",X"03",X"30",X"0C",X"7D",X"83",X"02",X"C9",X"F0",X"90",X"02",X"A9",
		X"00",X"B8",X"50",X"09",X"7D",X"83",X"02",X"C9",X"10",X"B0",X"02",X"A9",X"00",X"A8",X"BD",X"C3",
		X"02",X"18",X"7D",X"03",X"02",X"9D",X"03",X"02",X"BD",X"23",X"03",X"30",X"0C",X"7D",X"63",X"02",
		X"C9",X"F0",X"90",X"02",X"A0",X"00",X"B8",X"50",X"09",X"7D",X"63",X"02",X"C9",X"10",X"B0",X"02",
		X"A0",X"00",X"9D",X"63",X"02",X"BD",X"03",X"03",X"18",X"7D",X"43",X"02",X"9D",X"43",X"02",X"BD",
		X"63",X"03",X"30",X"0C",X"7D",X"A3",X"02",X"C9",X"F0",X"90",X"02",X"A0",X"00",X"B8",X"50",X"09",
		X"7D",X"A3",X"02",X"C9",X"10",X"B0",X"02",X"A0",X"00",X"9D",X"A3",X"02",X"98",X"9D",X"83",X"02",
		X"60",X"A9",X"FD",X"85",X"29",X"BD",X"C3",X"02",X"BC",X"23",X"03",X"20",X"5D",X"A7",X"9D",X"C3",
		X"02",X"98",X"9D",X"23",X"03",X"BD",X"E3",X"02",X"BC",X"43",X"03",X"20",X"5D",X"A7",X"9D",X"E3",
		X"02",X"98",X"9D",X"43",X"03",X"BD",X"03",X"03",X"BC",X"63",X"03",X"20",X"5D",X"A7",X"9D",X"03",
		X"03",X"98",X"9D",X"63",X"03",X"A5",X"29",X"D0",X"03",X"9D",X"83",X"02",X"60",X"84",X"2B",X"24",
		X"2B",X"30",X"0F",X"38",X"ED",X"88",X"A7",X"85",X"2A",X"A5",X"2B",X"E9",X"00",X"90",X"0F",X"B8",
		X"50",X"12",X"18",X"6D",X"88",X"A7",X"85",X"2A",X"A5",X"2B",X"69",X"00",X"90",X"06",X"E6",X"29",
		X"A9",X"00",X"85",X"2A",X"A8",X"A5",X"2A",X"60",X"20",X"A2",X"0F",X"A9",X"00",X"9D",X"83",X"02",
		X"CA",X"10",X"F8",X"A9",X"20",X"8D",X"0E",X"01",X"8D",X"0D",X"01",X"A9",X"04",X"85",X"01",X"A9",
		X"00",X"85",X"68",X"85",X"69",X"60",X"84",X"2A",X"38",X"E5",X"2A",X"85",X"2A",X"2C",X"11",X"01",
		X"30",X"09",X"29",X"0F",X"2C",X"BC",X"A7",X"F0",X"02",X"09",X"F8",X"60",X"08",X"A2",X"07",X"A9",
		X"00",X"9D",X"FE",X"03",X"CA",X"10",X"FA",X"A9",X"F0",X"8D",X"05",X"04",X"A9",X"FF",X"8D",X"15",
		X"01",X"60",X"AD",X"15",X"01",X"F0",X"59",X"A9",X"00",X"85",X"29",X"A2",X"07",X"86",X"37",X"A6",
		X"37",X"BD",X"FE",X"03",X"F0",X"18",X"38",X"E9",X"07",X"90",X"02",X"C9",X"10",X"B0",X"0C",X"AC",
		X"15",X"01",X"10",X"05",X"A9",X"F0",X"B8",X"50",X"02",X"A9",X"00",X"B8",X"50",X"20",X"AC",X"15",
		X"01",X"10",X"1B",X"8A",X"18",X"69",X"01",X"C9",X"08",X"90",X"02",X"A9",X"00",X"A8",X"B9",X"FE",
		X"03",X"F0",X"0B",X"C9",X"D5",X"B0",X"05",X"A9",X"F0",X"B8",X"50",X"02",X"A9",X"00",X"9D",X"FE",
		X"03",X"05",X"29",X"85",X"29",X"C6",X"37",X"10",X"B6",X"A5",X"29",X"D0",X"03",X"8D",X"15",X"01",
		X"60",X"A9",X"00",X"8D",X"AA",X"03",X"8D",X"25",X"01",X"60",X"A5",X"05",X"10",X"3E",X"AD",X"25",
		X"01",X"D0",X"23",X"AD",X"01",X"02",X"30",X"1B",X"A5",X"4E",X"29",X"08",X"F0",X"15",X"AD",X"AA",
		X"03",X"C9",X"02",X"B0",X"08",X"EE",X"AA",X"03",X"A9",X"01",X"8D",X"25",X"01",X"A5",X"4E",X"29",
		X"77",X"85",X"4E",X"B8",X"50",X"16",X"EE",X"25",X"01",X"AE",X"AA",X"03",X"AD",X"25",X"01",X"DD",
		X"83",X"A8",X"90",X"05",X"A9",X"00",X"8D",X"25",X"01",X"20",X"88",X"A8",X"A5",X"4E",X"29",X"7F",
		X"85",X"4E",X"60",X"00",X"13",X"05",X"00",X"00",X"AD",X"25",X"01",X"C9",X"03",X"90",X"14",X"29",
		X"01",X"D0",X"10",X"AC",X"1C",X"01",X"B9",X"DF",X"02",X"D0",X"09",X"88",X"10",X"F8",X"A9",X"00",
		X"8D",X"25",X"01",X"60",X"B9",X"8A",X"02",X"29",X"FC",X"99",X"8A",X"02",X"4C",X"98",X"A3",X"E1",
		X"24",X"26",X"28",X"2A",X"A9",X"01",X"85",X"72",X"20",X"6A",X"DF",X"A0",X"05",X"20",X"D1",X"B0",
		X"A5",X"05",X"30",X"26",X"A2",X"00",X"A5",X"03",X"29",X"20",X"D0",X"0C",X"A2",X"22",X"A5",X"06",
		X"F0",X"06",X"24",X"A2",X"30",X"02",X"A2",X"06",X"20",X"14",X"AB",X"20",X"0D",X"AB",X"AD",X"E4",
		X"31",X"8D",X"A6",X"2F",X"8D",X"A8",X"2F",X"20",X"A8",X"AA",X"A9",X"01",X"A0",X"00",X"20",X"7F",
		X"A9",X"24",X"05",X"30",X"09",X"A5",X"43",X"05",X"44",X"05",X"45",X"B8",X"50",X"02",X"A5",X"3E",
		X"F0",X"06",X"A9",X"01",X"A8",X"20",X"7F",X"A9",X"A5",X"00",X"C9",X"04",X"F0",X"35",X"A9",X"1D",
		X"85",X"3B",X"A9",X"07",X"85",X"3C",X"AE",X"E4",X"CD",X"20",X"D7",X"A9",X"A0",X"0A",X"A9",X"A7",
		X"59",X"CE",X"AA",X"88",X"10",X"FA",X"8D",X"6C",X"01",X"AE",X"E5",X"CD",X"A9",X"02",X"85",X"38",
		X"A4",X"38",X"B9",X"1B",X"06",X"0A",X"A8",X"B9",X"FA",X"31",X"9D",X"60",X"2F",X"E8",X"E8",X"C6",
		X"38",X"10",X"ED",X"A9",X"2F",X"A2",X"60",X"20",X"39",X"DF",X"AD",X"23",X"01",X"10",X"05",X"A2",
		X"36",X"20",X"14",X"AB",X"A5",X"00",X"C9",X"18",X"D0",X"22",X"A5",X"05",X"10",X"1E",X"A6",X"3D",
		X"BD",X"02",X"01",X"F0",X"0D",X"A2",X"30",X"20",X"14",X"AB",X"A4",X"3D",X"BE",X"02",X"01",X"20",
		X"C6",X"B0",X"A2",X"3A",X"20",X"14",X"AB",X"A2",X"38",X"20",X"14",X"AB",X"60",X"42",X"45",X"A6",
		X"00",X"E0",X"04",X"84",X"2B",X"C4",X"3D",X"D0",X"06",X"24",X"05",X"10",X"02",X"A9",X"00",X"09",
		X"70",X"BE",X"DE",X"CD",X"9D",X"60",X"2F",X"BE",X"E0",X"CD",X"B9",X"48",X"00",X"85",X"38",X"F0",
		X"06",X"C4",X"3D",X"D0",X"02",X"C6",X"38",X"A0",X"01",X"AD",X"84",X"32",X"C4",X"38",X"90",X"05",
		X"F0",X"03",X"AD",X"86",X"32",X"9D",X"60",X"2F",X"E8",X"E8",X"C8",X"C0",X"07",X"90",X"EA",X"A4",
		X"2B",X"A5",X"00",X"C9",X"04",X"D0",X"04",X"C4",X"3D",X"D0",X"30",X"BE",X"E2",X"CD",X"B9",X"7D",
		X"A9",X"85",X"3B",X"A9",X"00",X"85",X"3C",X"A0",X"02",X"84",X"2A",X"38",X"08",X"A0",X"00",X"B1",
		X"3B",X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"FC",X"A9",X"A5",X"2A",X"D0",X"01",X"18",X"A0",X"00",
		X"B1",X"3B",X"20",X"FC",X"A9",X"C6",X"3B",X"C6",X"2A",X"10",X"E1",X"60",X"29",X"0F",X"A8",X"F0",
		X"01",X"18",X"B0",X"01",X"C8",X"08",X"98",X"0A",X"A8",X"B9",X"E4",X"31",X"9D",X"60",X"2F",X"E8",
		X"E8",X"28",X"60",X"A6",X"3E",X"24",X"05",X"30",X"0A",X"A5",X"43",X"05",X"44",X"05",X"45",X"F0",
		X"02",X"A2",X"01",X"A9",X"60",X"85",X"74",X"A9",X"2F",X"85",X"75",X"BD",X"66",X"CE",X"A8",X"38",
		X"65",X"74",X"48",X"B9",X"E6",X"CD",X"91",X"74",X"88",X"D0",X"F8",X"B9",X"E6",X"CD",X"91",X"74",
		X"A5",X"05",X"10",X"10",X"A9",X"2F",X"85",X"75",X"A9",X"A6",X"85",X"74",X"A5",X"9F",X"18",X"69",
		X"01",X"20",X"77",X"AF",X"68",X"85",X"74",X"4C",X"09",X"DF",X"A2",X"08",X"20",X"14",X"AB",X"4C",
		X"69",X"AA",X"A9",X"30",X"A2",X"00",X"20",X"17",X"AB",X"20",X"92",X"AA",X"4C",X"E7",X"A8",X"20",
		X"B4",X"A8",X"A9",X"00",X"A2",X"06",X"4C",X"17",X"AB",X"A9",X"00",X"A2",X"32",X"20",X"17",X"AB",
		X"A5",X"03",X"29",X"1F",X"C9",X"10",X"B0",X"07",X"A9",X"E0",X"A2",X"22",X"20",X"17",X"AB",X"4C",
		X"B4",X"A8",X"A2",X"02",X"20",X"14",X"AB",X"A9",X"00",X"20",X"DD",X"B0",X"A6",X"3D",X"E8",X"86",
		X"61",X"A9",X"61",X"A0",X"01",X"4C",X"B1",X"DF",X"A5",X"09",X"29",X"03",X"AA",X"BD",X"B0",X"A8",
		X"AA",X"20",X"14",X"AB",X"CE",X"6E",X"01",X"A5",X"0A",X"29",X"01",X"F0",X"0E",X"A5",X"03",X"29",
		X"20",X"D0",X"08",X"A2",X"32",X"20",X"14",X"AB",X"B8",X"50",X"03",X"20",X"CA",X"AE",X"A2",X"2C",
		X"20",X"14",X"AB",X"A2",X"2E",X"20",X"14",X"AB",X"A5",X"06",X"C9",X"28",X"90",X"04",X"A9",X"28",
		X"85",X"06",X"20",X"77",X"AF",X"A5",X"17",X"F0",X"09",X"AD",X"F4",X"AA",X"AE",X"F3",X"AA",X"20",
		X"39",X"DF",X"60",X"5C",X"32",X"F8",X"85",X"29",X"A9",X"00",X"85",X"2C",X"A0",X"07",X"06",X"29",
		X"A5",X"2C",X"65",X"2C",X"85",X"2C",X"88",X"10",X"F5",X"D8",X"85",X"29",X"60",X"A9",X"20",X"A2",
		X"80",X"4C",X"57",X"DF",X"BD",X"22",X"D1",X"86",X"35",X"85",X"2B",X"A4",X"35",X"B1",X"AC",X"85",
		X"3B",X"C8",X"B1",X"AC",X"85",X"3C",X"E0",X"2C",X"D0",X"08",X"A5",X"74",X"85",X"B6",X"A5",X"75",
		X"85",X"B7",X"A0",X"00",X"B1",X"3B",X"85",X"2A",X"20",X"0D",X"AB",X"A9",X"00",X"85",X"73",X"A9",
		X"01",X"85",X"72",X"20",X"6A",X"DF",X"A5",X"2A",X"A6",X"2B",X"20",X"75",X"DF",X"A4",X"35",X"B1",
		X"AC",X"85",X"3B",X"C8",X"B1",X"AC",X"85",X"3C",X"A6",X"35",X"BD",X"21",X"D1",X"48",X"4A",X"4A",
		X"4A",X"4A",X"A8",X"20",X"D1",X"B0",X"68",X"29",X"0F",X"20",X"DD",X"B0",X"A0",X"01",X"A9",X"00",
		X"85",X"2A",X"B1",X"3B",X"85",X"2B",X"29",X"7F",X"C8",X"84",X"2C",X"AA",X"BD",X"E4",X"31",X"A4",
		X"2A",X"91",X"74",X"C8",X"BD",X"E5",X"31",X"91",X"74",X"C8",X"84",X"2A",X"A4",X"2C",X"24",X"2B",
		X"10",X"E0",X"A4",X"2A",X"88",X"4C",X"5F",X"DF",X"86",X"35",X"85",X"2A",X"A9",X"00",X"85",X"2B",
		X"F0",X"99",X"20",X"20",X"AC",X"AD",X"C9",X"01",X"29",X"03",X"F0",X"5B",X"20",X"20",X"AC",X"A9",
		X"08",X"8D",X"00",X"01",X"AD",X"1B",X"07",X"0D",X"1C",X"07",X"0D",X"1D",X"07",X"D0",X"03",X"20",
		X"36",X"AC",X"A2",X"17",X"AD",X"C9",X"01",X"29",X"01",X"D0",X"02",X"A2",X"0E",X"BD",X"08",X"AC",
		X"9D",X"06",X"06",X"CA",X"10",X"F7",X"A2",X"17",X"AD",X"C9",X"01",X"29",X"02",X"D0",X"02",X"A2",
		X"0E",X"A9",X"01",X"9D",X"06",X"07",X"CA",X"10",X"F8",X"AD",X"C9",X"01",X"29",X"03",X"F0",X"0F",
		X"A5",X"0A",X"29",X"F8",X"8D",X"1E",X"07",X"AD",X"6A",X"01",X"29",X"03",X"8D",X"1F",X"07",X"AD",
		X"C9",X"01",X"29",X"FC",X"8D",X"C9",X"01",X"60",X"07",X"04",X"01",X"0F",X"09",X"0C",X"0B",X"03",
		X"12",X"13",X"05",X"03",X"07",X"0F",X"0C",X"11",X"11",X"11",X"12",X"04",X"03",X"03",X"09",X"04",
		X"20",X"BB",X"D6",X"A5",X"0A",X"29",X"F8",X"CD",X"1E",X"07",X"D0",X"08",X"AD",X"6A",X"01",X"29",
		X"03",X"CD",X"1F",X"07",X"F0",X"08",X"AD",X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"60",X"A5",
		X"05",X"29",X"BF",X"85",X"05",X"A5",X"09",X"29",X"43",X"C9",X"40",X"D0",X"03",X"20",X"62",X"CA",
		X"20",X"FB",X"DD",X"A9",X"00",X"8D",X"01",X"06",X"A6",X"3E",X"F0",X"02",X"A2",X"03",X"B5",X"42",
		X"85",X"2C",X"B5",X"41",X"85",X"2D",X"B5",X"40",X"85",X"2E",X"8A",X"29",X"01",X"85",X"36",X"A9",
		X"00",X"85",X"2B",X"A9",X"1A",X"85",X"2A",X"85",X"29",X"A9",X"00",X"8D",X"05",X"06",X"A0",X"FD",
		X"B9",X"20",X"06",X"C5",X"2C",X"D0",X"14",X"B9",X"1F",X"06",X"C5",X"2D",X"D0",X"0D",X"C0",X"52",
		X"90",X"08",X"B9",X"1E",X"06",X"C5",X"2E",X"B8",X"50",X"01",X"38",X"B0",X"4F",X"C0",X"E8",X"90",
		X"1E",X"A5",X"29",X"BE",X"1E",X"05",X"99",X"1E",X"05",X"86",X"29",X"A5",X"2A",X"BE",X"1F",X"05",
		X"99",X"1F",X"05",X"86",X"2A",X"A5",X"2B",X"BE",X"20",X"05",X"99",X"20",X"05",X"86",X"2B",X"A5",
		X"2D",X"BE",X"1F",X"06",X"99",X"1F",X"06",X"86",X"2D",X"A5",X"2C",X"BE",X"20",X"06",X"99",X"20",
		X"06",X"86",X"2C",X"C0",X"52",X"90",X"0A",X"A5",X"2E",X"BE",X"1E",X"06",X"99",X"1E",X"06",X"86",
		X"2E",X"C0",X"55",X"90",X"01",X"88",X"88",X"88",X"D0",X"B3",X"A0",X"02",X"EE",X"05",X"06",X"C0",
		X"55",X"90",X"01",X"88",X"88",X"88",X"D0",X"88",X"A6",X"36",X"AD",X"05",X"06",X"9D",X"00",X"06",
		X"CA",X"30",X"03",X"4C",X"5E",X"AC",X"AD",X"01",X"06",X"CD",X"00",X"06",X"90",X"07",X"C9",X"63",
		X"B0",X"03",X"EE",X"01",X"06",X"A5",X"3D",X"49",X"01",X"0A",X"0A",X"05",X"3D",X"69",X"05",X"8D",
		X"03",X"06",X"A0",X"14",X"AD",X"03",X"06",X"F0",X"42",X"29",X"03",X"85",X"3D",X"C6",X"3D",X"4E",
		X"03",X"06",X"4E",X"03",X"06",X"A6",X"3D",X"BD",X"00",X"06",X"F0",X"2C",X"C9",X"09",X"B0",X"28",
		X"0A",X"18",X"7D",X"00",X"06",X"49",X"FF",X"38",X"E9",X"E5",X"8D",X"02",X"06",X"20",X"48",X"CA",
		X"A9",X"60",X"8D",X"05",X"06",X"A9",X"00",X"85",X"4E",X"85",X"50",X"A9",X"02",X"8D",X"04",X"06",
		X"20",X"89",X"A7",X"A0",X"24",X"84",X"00",X"60",X"4C",X"22",X"AD",X"84",X"00",X"60",X"A9",X"06",
		X"85",X"01",X"A5",X"03",X"29",X"1F",X"D0",X"0A",X"CE",X"05",X"06",X"D0",X"05",X"A0",X"14",X"84",
		X"00",X"60",X"AE",X"02",X"06",X"BD",X"06",X"06",X"20",X"CE",X"AD",X"A8",X"10",X"05",X"A9",X"1A",
		X"B8",X"50",X"06",X"C9",X"1B",X"90",X"02",X"A9",X"00",X"AE",X"02",X"06",X"9D",X"06",X"06",X"A5",
		X"4E",X"29",X"18",X"A8",X"A5",X"4E",X"29",X"67",X"85",X"4E",X"98",X"F0",X"20",X"CE",X"02",X"06",
		X"CE",X"04",X"06",X"10",X"12",X"A6",X"3D",X"BD",X"00",X"06",X"C9",X"04",X"B0",X"03",X"20",X"F7",
		X"DD",X"20",X"22",X"AD",X"B8",X"50",X"06",X"CA",X"A9",X"00",X"9D",X"06",X"06",X"60",X"48",X"A5",
		X"50",X"0A",X"0A",X"0A",X"18",X"65",X"51",X"85",X"51",X"68",X"A4",X"50",X"30",X"05",X"69",X"00",
		X"B8",X"50",X"02",X"69",X"FF",X"A0",X"00",X"84",X"50",X"60",X"20",X"B4",X"A8",X"A9",X"C0",X"A2",
		X"02",X"20",X"17",X"AB",X"CE",X"6E",X"01",X"20",X"97",X"AA",X"A2",X"0A",X"20",X"14",X"AB",X"A9",
		X"A6",X"A2",X"0C",X"20",X"17",X"AB",X"A9",X"9C",X"A2",X"0E",X"20",X"17",X"AB",X"A2",X"2C",X"20",
		X"14",X"AB",X"AD",X"02",X"06",X"38",X"ED",X"04",X"06",X"4C",X"4E",X"AE",X"20",X"B4",X"A8",X"78",
		X"AD",X"CA",X"60",X"AC",X"CA",X"60",X"84",X"29",X"4A",X"4A",X"4A",X"4A",X"45",X"29",X"85",X"29",
		X"AD",X"DA",X"60",X"AC",X"DA",X"60",X"58",X"45",X"29",X"29",X"F0",X"45",X"29",X"85",X"29",X"98",
		X"0A",X"0A",X"0A",X"0A",X"45",X"29",X"8D",X"1F",X"01",X"20",X"26",X"AF",X"A9",X"FF",X"85",X"63",
		X"A2",X"10",X"20",X"14",X"AB",X"A9",X"01",X"85",X"61",X"20",X"DD",X"B0",X"A9",X"28",X"85",X"2C",
		X"A2",X"15",X"86",X"37",X"20",X"0D",X"AB",X"A9",X"00",X"85",X"73",X"A5",X"2C",X"AA",X"38",X"E9",
		X"0A",X"85",X"2C",X"A9",X"D0",X"20",X"75",X"DF",X"A0",X"07",X"A5",X"63",X"C5",X"37",X"D0",X"02",
		X"A0",X"00",X"20",X"D1",X"B0",X"A9",X"61",X"A0",X"01",X"20",X"B1",X"DF",X"A9",X"A0",X"20",X"6A",
		X"B5",X"A9",X"00",X"85",X"73",X"AA",X"A9",X"08",X"20",X"75",X"DF",X"E6",X"61",X"A5",X"37",X"20",
		X"F8",X"AE",X"A2",X"00",X"A9",X"08",X"20",X"75",X"DF",X"A6",X"37",X"BD",X"06",X"07",X"85",X"56",
		X"BD",X"07",X"07",X"85",X"57",X"BD",X"08",X"07",X"85",X"58",X"A9",X"56",X"A0",X"03",X"20",X"B1",
		X"DF",X"C6",X"37",X"C6",X"37",X"C6",X"37",X"10",X"9B",X"60",X"AD",X"56",X"01",X"F0",X"14",X"85",
		X"58",X"A2",X"34",X"20",X"14",X"AB",X"A9",X"00",X"85",X"56",X"85",X"57",X"A9",X"56",X"A0",X"03",
		X"20",X"B1",X"DF",X"18",X"A0",X"10",X"A9",X"85",X"79",X"75",X"D5",X"88",X"10",X"FA",X"85",X"B5",
		X"60",X"AD",X"02",X"06",X"38",X"ED",X"04",X"06",X"18",X"69",X"02",X"85",X"38",X"A0",X"00",X"A9",
		X"02",X"85",X"39",X"A6",X"38",X"BD",X"06",X"06",X"C9",X"1E",X"90",X"02",X"A9",X"1A",X"0A",X"AA",
		X"BD",X"FA",X"31",X"91",X"74",X"C8",X"BD",X"FB",X"31",X"91",X"74",X"C8",X"C6",X"38",X"C6",X"39",
		X"10",X"E1",X"88",X"4C",X"5F",X"DF",X"AD",X"00",X"06",X"0D",X"01",X"06",X"F0",X"40",X"A2",X"12",
		X"20",X"14",X"AB",X"A9",X"63",X"20",X"71",X"AF",X"A2",X"00",X"20",X"3F",X"AF",X"A2",X"01",X"BD",
		X"00",X"06",X"F0",X"2A",X"48",X"86",X"2E",X"A0",X"03",X"20",X"D1",X"B0",X"20",X"0D",X"AB",X"A9",
		X"D0",X"A4",X"2E",X"BE",X"6F",X"AF",X"20",X"75",X"DF",X"68",X"20",X"71",X"AF",X"A9",X"A0",X"20",
		X"6A",X"B5",X"A9",X"10",X"A2",X"04",X"20",X"98",X"AB",X"A6",X"2E",X"20",X"9E",X"AA",X"60",X"C0",
		X"B0",X"C9",X"63",X"90",X"02",X"A9",X"63",X"20",X"F5",X"AA",X"A9",X"29",X"A0",X"01",X"4C",X"B1",
		X"DF",X"20",X"48",X"CA",X"CE",X"6E",X"01",X"A0",X"03",X"20",X"D1",X"B0",X"A9",X"01",X"85",X"72",
		X"20",X"6A",X"DF",X"A2",X"2C",X"A9",X"60",X"20",X"17",X"AB",X"20",X"92",X"AA",X"A2",X"07",X"86",
		X"37",X"A4",X"37",X"BE",X"9B",X"B0",X"20",X"14",X"AB",X"C6",X"37",X"10",X"F4",X"AD",X"00",X"02",
		X"38",X"E5",X"7B",X"10",X"07",X"C6",X"7B",X"C6",X"7C",X"B8",X"50",X"25",X"D0",X"0D",X"C6",X"7C",
		X"C6",X"7B",X"10",X"04",X"E6",X"7B",X"E6",X"7C",X"B8",X"50",X"16",X"A5",X"7C",X"CD",X"27",X"01",
		X"F0",X"02",X"B0",X"0D",X"38",X"ED",X"00",X"02",X"D0",X"01",X"18",X"B0",X"04",X"E6",X"7B",X"E6",
		X"7C",X"A5",X"7C",X"85",X"3A",X"A2",X"04",X"86",X"37",X"A0",X"05",X"20",X"D1",X"B0",X"A9",X"00",
		X"85",X"73",X"20",X"0D",X"AB",X"A2",X"D8",X"A4",X"37",X"B9",X"96",X"B0",X"18",X"69",X"F8",X"20",
		X"75",X"DF",X"A6",X"3A",X"BC",X"FE",X"91",X"C0",X"63",X"B0",X"37",X"C8",X"98",X"20",X"77",X"AF",
		X"A0",X"03",X"20",X"D1",X"B0",X"20",X"0D",X"AB",X"A2",X"BA",X"A4",X"37",X"B9",X"96",X"B0",X"18",
		X"69",X"EC",X"20",X"75",X"DF",X"A6",X"3A",X"20",X"C6",X"B0",X"20",X"0D",X"AB",X"A2",X"CC",X"A4",
		X"37",X"B9",X"96",X"B0",X"18",X"69",X"00",X"20",X"75",X"DF",X"A6",X"3A",X"BD",X"FE",X"91",X"20",
		X"E1",X"C4",X"C6",X"3A",X"C6",X"37",X"10",X"A1",X"A9",X"00",X"85",X"73",X"20",X"0D",X"AB",X"A2",
		X"1C",X"20",X"14",X"AB",X"A9",X"04",X"A0",X"01",X"20",X"B1",X"DF",X"A0",X"00",X"20",X"D1",X"B0",
		X"20",X"0D",X"AB",X"A2",X"B8",X"20",X"AB",X"B0",X"38",X"E5",X"7B",X"A8",X"B9",X"96",X"B0",X"38",
		X"E9",X"16",X"20",X"75",X"DF",X"A9",X"E0",X"85",X"73",X"A2",X"00",X"86",X"38",X"A0",X"03",X"84",
		X"37",X"A4",X"38",X"B9",X"A3",X"B0",X"AA",X"C8",X"B9",X"A3",X"B0",X"C8",X"84",X"38",X"20",X"75",
		X"DF",X"C6",X"37",X"10",X"EC",X"60",X"BE",X"E3",X"09",X"30",X"58",X"14",X"0C",X"0E",X"16",X"18",
		X"1E",X"20",X"1A",X"00",X"26",X"28",X"00",X"00",X"DA",X"D8",X"00",X"AD",X"00",X"02",X"20",X"CE",
		X"AD",X"A8",X"10",X"05",X"A9",X"00",X"B8",X"50",X"08",X"CD",X"27",X"01",X"90",X"03",X"AD",X"27",
		X"01",X"8D",X"00",X"02",X"A8",X"60",X"8A",X"20",X"B5",X"91",X"A9",X"29",X"A0",X"03",X"4C",X"B1",
		X"DF",X"C4",X"9E",X"F0",X"07",X"84",X"9E",X"A9",X"08",X"4C",X"4C",X"DF",X"60",X"C5",X"72",X"F0",
		X"05",X"85",X"72",X"4C",X"6A",X"DF",X"60",X"A9",X"0A",X"85",X"00",X"A9",X"00",X"85",X"02",X"A9",
		X"DF",X"85",X"04",X"A9",X"12",X"85",X"01",X"A9",X"19",X"8D",X"4E",X"01",X"A9",X"18",X"8D",X"4D",
		X"01",X"60",X"A9",X"34",X"A2",X"AA",X"20",X"5A",X"B1",X"AD",X"4E",X"01",X"C9",X"A0",X"B0",X"05",
		X"69",X"14",X"8D",X"4E",X"01",X"C9",X"50",X"90",X"17",X"AD",X"4D",X"01",X"18",X"69",X"08",X"8D",
		X"4D",X"01",X"CD",X"4E",X"01",X"90",X"09",X"A9",X"A0",X"8D",X"4D",X"01",X"A9",X"14",X"85",X"01",
		X"60",X"A9",X"3F",X"A2",X"4E",X"20",X"5A",X"B1",X"AD",X"4D",X"01",X"C9",X"30",X"90",X"05",X"E9",
		X"01",X"8D",X"4D",X"01",X"C9",X"80",X"B0",X"11",X"AD",X"4E",X"01",X"38",X"E9",X"01",X"CD",X"4D",
		X"01",X"B0",X"03",X"AD",X"4D",X"01",X"8D",X"4E",X"01",X"60",X"85",X"57",X"86",X"56",X"AD",X"4D",
		X"01",X"85",X"37",X"CE",X"6E",X"01",X"A5",X"37",X"0A",X"0A",X"29",X"7F",X"A8",X"A5",X"37",X"4A",
		X"4A",X"4A",X"4A",X"4A",X"20",X"6C",X"DF",X"A5",X"37",X"CD",X"4D",X"01",X"D0",X"05",X"A9",X"00",
		X"B8",X"50",X"0C",X"4A",X"4A",X"4A",X"EA",X"29",X"07",X"C9",X"07",X"D0",X"02",X"A9",X"03",X"A8",
		X"A9",X"68",X"20",X"4C",X"DF",X"A5",X"57",X"A6",X"56",X"20",X"39",X"DF",X"A5",X"37",X"18",X"69",
		X"02",X"85",X"37",X"CD",X"4E",X"01",X"90",X"BE",X"A2",X"2C",X"A9",X"D0",X"20",X"17",X"AB",X"A9",
		X"3F",X"A2",X"F2",X"4C",X"39",X"DF",X"20",X"C3",X"C1",X"AD",X"00",X"20",X"CD",X"C6",X"CE",X"D0",
		X"06",X"AD",X"33",X"01",X"D0",X"01",X"60",X"A5",X"01",X"C9",X"00",X"F0",X"3C",X"A9",X"00",X"20",
		X"BE",X"B2",X"20",X"32",X"B3",X"B0",X"1E",X"20",X"0D",X"B2",X"AD",X"6E",X"01",X"F0",X"16",X"A0",
		X"27",X"A9",X"0E",X"38",X"F1",X"B6",X"88",X"10",X"FB",X"A8",X"F0",X"02",X"49",X"E5",X"F0",X"02",
		X"49",X"29",X"8D",X"55",X"04",X"A9",X"00",X"20",X"FE",X"B2",X"AD",X"C4",X"CE",X"8D",X"00",X"20",
		X"AD",X"C5",X"CE",X"8D",X"01",X"20",X"B8",X"50",X"03",X"4C",X"30",X"B2",X"60",X"A6",X"01",X"BD",
		X"19",X"B2",X"48",X"BD",X"18",X"B2",X"48",X"60",X"2F",X"B2",X"03",X"D8",X"B9",X"B8",X"E9",X"AD",
		X"80",X"AF",X"1B",X"AE",X"61",X"AA",X"59",X"AA",X"6E",X"AA",X"01",X"B1",X"30",X"B1",X"78",X"AA",
		X"A9",X"07",X"20",X"BE",X"B2",X"20",X"86",X"B5",X"A9",X"07",X"20",X"FE",X"B2",X"A9",X"04",X"20",
		X"BE",X"B2",X"20",X"5B",X"B7",X"A9",X"04",X"20",X"FE",X"B2",X"A9",X"03",X"20",X"BE",X"B2",X"20",
		X"AD",X"B5",X"A9",X"03",X"20",X"FE",X"B2",X"A9",X"06",X"20",X"BE",X"B2",X"20",X"9A",X"B7",X"A9",
		X"06",X"20",X"FE",X"B2",X"A9",X"05",X"20",X"BE",X"B2",X"20",X"98",X"B4",X"A9",X"05",X"20",X"FE",
		X"B2",X"A9",X"00",X"20",X"BE",X"B2",X"20",X"B4",X"A8",X"A5",X"05",X"30",X"0D",X"A9",X"F2",X"18",
		X"A0",X"27",X"71",X"B6",X"88",X"10",X"FB",X"8D",X"1B",X"01",X"A9",X"00",X"20",X"FE",X"B2",X"20",
		X"67",X"B3",X"A9",X"01",X"20",X"BE",X"B2",X"20",X"C2",X"C5",X"A9",X"01",X"20",X"FE",X"B2",X"A9",
		X"08",X"20",X"BE",X"B2",X"20",X"4D",X"C5",X"A9",X"08",X"20",X"FE",X"B2",X"A9",X"00",X"8D",X"14",
		X"01",X"AD",X"C2",X"CE",X"8D",X"00",X"20",X"AD",X"C3",X"CE",X"8D",X"01",X"20",X"60",X"AA",X"0A",
		X"A8",X"BD",X"15",X"04",X"D0",X"09",X"BE",X"7A",X"CE",X"B9",X"7B",X"CE",X"B8",X"50",X"06",X"BE",
		X"68",X"CE",X"B9",X"69",X"CE",X"86",X"74",X"85",X"75",X"A9",X"00",X"85",X"A9",X"60",X"AA",X"0A",
		X"A8",X"BD",X"15",X"04",X"D0",X"09",X"BE",X"68",X"CE",X"B9",X"69",X"CE",X"B8",X"50",X"06",X"BE",
		X"7A",X"CE",X"B9",X"7B",X"CE",X"86",X"3B",X"85",X"3C",X"A9",X"00",X"85",X"A9",X"60",X"48",X"20",
		X"09",X"DF",X"68",X"AA",X"0A",X"A8",X"B9",X"8C",X"CE",X"85",X"3B",X"B9",X"8D",X"CE",X"85",X"3C",
		X"BD",X"15",X"04",X"49",X"01",X"9D",X"15",X"04",X"D0",X"09",X"B9",X"9E",X"CE",X"BE",X"9F",X"CE",
		X"B8",X"50",X"06",X"B9",X"B0",X"CE",X"BE",X"B1",X"CE",X"A0",X"00",X"91",X"3B",X"8A",X"C8",X"91",
		X"3B",X"60",X"AD",X"C4",X"CE",X"CD",X"00",X"20",X"F0",X"05",X"8D",X"00",X"20",X"38",X"60",X"AD",
		X"15",X"04",X"D0",X"05",X"A2",X"02",X"B8",X"50",X"02",X"A2",X"08",X"BD",X"9E",X"CE",X"A0",X"00",
		X"8C",X"6E",X"01",X"91",X"74",X"C8",X"BD",X"9F",X"CE",X"91",X"74",X"BD",X"68",X"CE",X"85",X"74",
		X"BD",X"69",X"CE",X"85",X"75",X"18",X"60",X"AD",X"14",X"01",X"F0",X"0D",X"A9",X"02",X"20",X"BE",
		X"B2",X"20",X"0D",X"C3",X"A9",X"02",X"20",X"FE",X"B2",X"A9",X"02",X"20",X"DE",X"B2",X"A9",X"00",
		X"A2",X"0F",X"9D",X"25",X"04",X"CA",X"10",X"FA",X"AD",X"06",X"01",X"30",X"49",X"AE",X"1C",X"01",
		X"BD",X"DF",X"02",X"F0",X"3E",X"A0",X"00",X"BD",X"83",X"02",X"29",X"07",X"C9",X"01",X"D0",X"33",
		X"C8",X"84",X"29",X"BD",X"83",X"02",X"29",X"80",X"D0",X"1C",X"AD",X"48",X"01",X"30",X"0C",X"BD",
		X"DF",X"02",X"CD",X"57",X"01",X"B0",X"04",X"E6",X"29",X"E6",X"29",X"A5",X"29",X"BC",X"CC",X"02",
		X"19",X"25",X"04",X"99",X"25",X"04",X"BC",X"B9",X"02",X"A5",X"29",X"09",X"80",X"19",X"25",X"04",
		X"99",X"25",X"04",X"CA",X"10",X"BA",X"A9",X"06",X"AC",X"25",X"01",X"F0",X"0C",X"30",X"0A",X"A5",
		X"03",X"29",X"07",X"C9",X"07",X"D0",X"02",X"A9",X"01",X"85",X"29",X"A0",X"FF",X"A2",X"FF",X"86",
		X"2C",X"AD",X"02",X"02",X"F0",X"0B",X"AD",X"01",X"02",X"30",X"06",X"AE",X"00",X"02",X"AC",X"01",
		X"02",X"86",X"2A",X"84",X"2B",X"AD",X"24",X"01",X"30",X"08",X"29",X"0E",X"4A",X"85",X"2C",X"CE",
		X"24",X"01",X"A2",X"0F",X"A0",X"06",X"BD",X"25",X"04",X"F0",X"0C",X"29",X"02",X"F0",X"05",X"A5",
		X"03",X"29",X"01",X"A8",X"B8",X"50",X"24",X"E4",X"2A",X"F0",X"02",X"E4",X"2B",X"D0",X"05",X"A0",
		X"01",X"B8",X"50",X"17",X"AD",X"24",X"01",X"30",X"10",X"8A",X"18",X"65",X"2C",X"29",X"07",X"C9",
		X"07",X"D0",X"02",X"A9",X"03",X"A8",X"B8",X"50",X"02",X"A4",X"29",X"98",X"BC",X"76",X"B4",X"91",
		X"3B",X"CA",X"10",X"C0",X"A2",X"0F",X"2C",X"11",X"01",X"10",X"01",X"CA",X"A0",X"C0",X"BD",X"25",
		X"04",X"10",X"02",X"A0",X"00",X"84",X"58",X"BC",X"87",X"B4",X"B1",X"B0",X"29",X"1F",X"05",X"58",
		X"91",X"B0",X"CA",X"10",X"E7",X"60",X"A8",X"9C",X"92",X"86",X"7C",X"70",X"66",X"5A",X"50",X"44",
		X"3A",X"2E",X"24",X"18",X"0E",X"02",X"B2",X"3B",X"37",X"33",X"2F",X"2B",X"27",X"23",X"1F",X"1B",
		X"17",X"13",X"0F",X"0B",X"07",X"03",X"3F",X"1D",X"A0",X"0C",X"84",X"9E",X"A9",X"08",X"20",X"4C",
		X"DF",X"A2",X"66",X"20",X"65",X"C7",X"A9",X"12",X"85",X"56",X"A2",X"3F",X"86",X"37",X"A0",X"00",
		X"A6",X"37",X"BD",X"43",X"02",X"D0",X"03",X"4C",X"49",X"B5",X"C9",X"50",X"90",X"02",X"C6",X"37",
		X"48",X"29",X"3F",X"91",X"74",X"68",X"2A",X"2A",X"2A",X"29",X"03",X"18",X"69",X"01",X"09",X"70",
		X"C8",X"91",X"74",X"C8",X"BD",X"03",X"02",X"AA",X"BD",X"8A",X"03",X"38",X"E5",X"68",X"85",X"63",
		X"91",X"74",X"C8",X"BD",X"7A",X"03",X"E5",X"69",X"85",X"64",X"29",X"1F",X"91",X"74",X"C8",X"BD",
		X"6A",X"03",X"85",X"61",X"91",X"74",X"C8",X"BD",X"5A",X"03",X"85",X"62",X"29",X"1F",X"91",X"74",
		X"C8",X"A9",X"00",X"91",X"74",X"C8",X"91",X"74",X"C8",X"91",X"74",X"A9",X"A0",X"C8",X"91",X"74",
		X"C8",X"A5",X"63",X"49",X"FF",X"18",X"69",X"01",X"91",X"74",X"C8",X"A5",X"64",X"49",X"FF",X"69",
		X"00",X"29",X"1F",X"91",X"74",X"C8",X"A5",X"61",X"49",X"FF",X"18",X"69",X"01",X"91",X"74",X"C8",
		X"A5",X"62",X"49",X"FF",X"69",X"00",X"29",X"1F",X"91",X"74",X"C8",X"C0",X"F0",X"90",X"06",X"88",
		X"20",X"5F",X"DF",X"A0",X"00",X"C6",X"56",X"30",X"07",X"C6",X"37",X"30",X"03",X"4C",X"B0",X"B4",
		X"98",X"F0",X"04",X"88",X"20",X"5F",X"DF",X"A5",X"B5",X"F0",X"0A",X"A5",X"46",X"C9",X"0A",X"90",
		X"04",X"A9",X"7A",X"85",X"53",X"A9",X"01",X"4C",X"6A",X"DF",X"48",X"A0",X"00",X"98",X"91",X"74",
		X"C8",X"91",X"74",X"C8",X"91",X"74",X"C8",X"68",X"91",X"74",X"A9",X"04",X"18",X"65",X"74",X"85",
		X"74",X"90",X"02",X"E6",X"75",X"60",X"A9",X"01",X"85",X"9E",X"AD",X"02",X"02",X"F0",X"1D",X"C9",
		X"F0",X"B0",X"19",X"85",X"57",X"85",X"2F",X"AD",X"01",X"02",X"C9",X"81",X"F0",X"0E",X"AC",X"00",
		X"02",X"A5",X"51",X"4A",X"29",X"07",X"18",X"69",X"01",X"20",X"A0",X"BD",X"60",X"AD",X"06",X"01",
		X"30",X"24",X"A2",X"06",X"86",X"37",X"A6",X"37",X"BD",X"DF",X"02",X"F0",X"15",X"85",X"57",X"BD",
		X"83",X"02",X"29",X"18",X"4A",X"4A",X"4A",X"85",X"55",X"BD",X"83",X"02",X"29",X"07",X"0A",X"20",
		X"D7",X"B5",X"C6",X"37",X"10",X"E0",X"60",X"A8",X"B9",X"E2",X"B5",X"48",X"B9",X"E1",X"B5",X"48",
		X"60",X"EA",X"B5",X"1A",X"B7",X"0E",X"B6",X"21",X"B6",X"9A",X"B6",X"A9",X"03",X"85",X"9E",X"BD",
		X"83",X"02",X"30",X"0E",X"BC",X"B9",X"02",X"A6",X"55",X"BD",X"0B",X"B6",X"20",X"A0",X"BD",X"B8",
		X"50",X"08",X"20",X"34",X"B6",X"A0",X"00",X"20",X"CB",X"BD",X"60",X"00",X"00",X"00",X"00",X"BD",
		X"8A",X"02",X"29",X"03",X"A8",X"B9",X"1E",X"B6",X"BC",X"B9",X"02",X"4C",X"FD",X"BC",X"1A",X"1A",
		X"4A",X"4C",X"BC",X"B9",X"02",X"A5",X"03",X"29",X"03",X"0A",X"18",X"69",X"12",X"4C",X"FD",X"BC",
		X"12",X"14",X"16",X"18",X"A5",X"57",X"85",X"2F",X"BC",X"B9",X"02",X"B9",X"CE",X"03",X"85",X"56",
		X"B9",X"DE",X"03",X"85",X"58",X"BD",X"CC",X"02",X"29",X"0F",X"A8",X"A5",X"56",X"49",X"80",X"18",
		X"79",X"8B",X"B6",X"50",X"09",X"10",X"05",X"A9",X"7F",X"B8",X"50",X"02",X"A9",X"80",X"49",X"80",
		X"85",X"2E",X"A5",X"58",X"49",X"80",X"18",X"79",X"87",X"B6",X"50",X"09",X"10",X"05",X"A9",X"7F",
		X"B8",X"50",X"02",X"A9",X"80",X"49",X"80",X"85",X"30",X"AC",X"12",X"01",X"B9",X"DC",X"BC",X"85",
		X"59",X"B9",X"EC",X"BC",X"85",X"5A",X"60",X"00",X"10",X"1F",X"28",X"2C",X"28",X"1F",X"10",X"00",
		X"F0",X"E1",X"D8",X"D4",X"D8",X"E1",X"F0",X"00",X"10",X"1F",X"28",X"BD",X"DF",X"02",X"85",X"57",
		X"BC",X"B9",X"02",X"B9",X"CE",X"03",X"85",X"56",X"B9",X"DE",X"03",X"85",X"58",X"BD",X"CC",X"02",
		X"10",X"23",X"98",X"18",X"69",X"01",X"29",X"0F",X"A8",X"B9",X"CE",X"03",X"38",X"E5",X"56",X"20",
		X"FA",X"B6",X"18",X"65",X"56",X"85",X"56",X"B9",X"DE",X"03",X"38",X"E5",X"58",X"20",X"FA",X"B6",
		X"18",X"65",X"58",X"85",X"58",X"20",X"98",X"C0",X"A2",X"61",X"20",X"65",X"C7",X"A9",X"00",X"85",
		X"A9",X"20",X"3E",X"BD",X"84",X"A9",X"A5",X"03",X"29",X"03",X"0A",X"18",X"69",X"4E",X"A8",X"BE",
		X"C9",X"CE",X"B9",X"C8",X"CE",X"A4",X"A9",X"4C",X"59",X"DF",X"85",X"29",X"BD",X"CC",X"02",X"29",
		X"07",X"85",X"2C",X"86",X"2B",X"A2",X"02",X"A9",X"00",X"46",X"2C",X"90",X"03",X"18",X"65",X"29",
		X"0A",X"08",X"6A",X"28",X"6A",X"CA",X"10",X"F1",X"A6",X"2B",X"60",X"A9",X"04",X"AC",X"48",X"01",
		X"30",X"02",X"A9",X"00",X"85",X"9E",X"AD",X"48",X"01",X"18",X"69",X"40",X"4A",X"4A",X"4A",X"4A",
		X"C9",X"05",X"90",X"02",X"A9",X"00",X"A8",X"B9",X"55",X"B7",X"85",X"29",X"BD",X"83",X"02",X"30",
		X"0B",X"BC",X"B9",X"02",X"A5",X"29",X"20",X"A0",X"BD",X"B8",X"50",X"08",X"20",X"34",X"B6",X"A4",
		X"29",X"20",X"CB",X"BD",X"60",X"0D",X"0C",X"0B",X"0A",X"09",X"09",X"A2",X"0B",X"86",X"37",X"A6",
		X"37",X"BD",X"D3",X"02",X"F0",X"1B",X"85",X"57",X"85",X"2F",X"E0",X"08",X"BC",X"AD",X"02",X"B0",
		X"05",X"A9",X"08",X"B8",X"50",X"08",X"A5",X"03",X"0A",X"29",X"06",X"18",X"69",X"20",X"20",X"FD",
		X"BC",X"C6",X"37",X"10",X"DA",X"A0",X"04",X"AD",X"35",X"01",X"C9",X"06",X"90",X"08",X"A0",X"0B",
		X"C9",X"08",X"90",X"02",X"A0",X"0C",X"8C",X"08",X"08",X"60",X"A0",X"00",X"84",X"9E",X"A2",X"07",
		X"86",X"37",X"A6",X"37",X"BD",X"0A",X"03",X"F0",X"29",X"85",X"57",X"BD",X"FA",X"02",X"85",X"29",
		X"BC",X"02",X"03",X"C0",X"01",X"D0",X"06",X"20",X"EB",X"B7",X"B8",X"50",X"15",X"BD",X"12",X"03",
		X"4A",X"29",X"FE",X"C0",X"02",X"90",X"02",X"A9",X"00",X"18",X"79",X"E5",X"B7",X"A4",X"29",X"20",
		X"FD",X"BC",X"C6",X"37",X"10",X"CC",X"AD",X"20",X"07",X"F0",X"09",X"A5",X"9F",X"C9",X"0D",X"90",
		X"03",X"8D",X"FF",X"01",X"60",X"00",X"00",X"5A",X"58",X"56",X"1C",X"A4",X"29",X"B9",X"35",X"04",
		X"85",X"56",X"B9",X"45",X"04",X"85",X"58",X"20",X"98",X"C0",X"A2",X"61",X"20",X"65",X"C7",X"AE",
		X"3B",X"01",X"CE",X"3C",X"01",X"D0",X"0A",X"E8",X"8E",X"3B",X"01",X"BD",X"2A",X"B8",X"8D",X"3C",
		X"01",X"BC",X"3D",X"B8",X"30",X"03",X"20",X"4E",X"B8",X"AD",X"3B",X"01",X"0A",X"18",X"69",X"28",
		X"A8",X"BE",X"C9",X"CE",X"B9",X"C8",X"CE",X"4C",X"57",X"DF",X"02",X"02",X"02",X"02",X"02",X"04",
		X"03",X"02",X"01",X"20",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"3B",X"B8",X"00",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"04",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B9",X"58",
		X"B8",X"48",X"B9",X"57",X"B8",X"48",X"60",X"5E",X"B8",X"74",X"B8",X"87",X"B8",X"95",X"B8",X"A9",
		X"0C",X"8D",X"0B",X"08",X"85",X"24",X"A9",X"04",X"8D",X"0A",X"08",X"85",X"23",X"A9",X"00",X"85",
		X"22",X"8D",X"09",X"08",X"60",X"A4",X"22",X"A2",X"02",X"B5",X"22",X"48",X"94",X"22",X"98",X"9D",
		X"09",X"08",X"68",X"A8",X"CA",X"10",X"F2",X"60",X"20",X"96",X"C1",X"A9",X"7F",X"8D",X"39",X"01",
		X"A9",X"04",X"8D",X"3A",X"01",X"60",X"AD",X"39",X"01",X"8D",X"FC",X"2F",X"AD",X"3A",X"01",X"09",
		X"70",X"8D",X"FD",X"2F",X"A9",X"C0",X"8D",X"FF",X"2F",X"AD",X"39",X"01",X"38",X"E9",X"20",X"10",
		X"05",X"29",X"7F",X"CE",X"3A",X"01",X"8D",X"39",X"01",X"60",X"A9",X"3F",X"A2",X"F2",X"20",X"39",
		X"DF",X"A9",X"00",X"85",X"6A",X"85",X"6B",X"85",X"6C",X"85",X"6D",X"8D",X"02",X"02",X"85",X"68",
		X"85",X"69",X"A9",X"E0",X"85",X"5F",X"A9",X"FF",X"85",X"5B",X"20",X"67",X"B9",X"85",X"77",X"86",
		X"76",X"A2",X"0F",X"86",X"37",X"A6",X"37",X"BD",X"83",X"02",X"F0",X"49",X"85",X"57",X"BD",X"63",
		X"02",X"85",X"56",X"BD",X"A3",X"02",X"85",X"58",X"20",X"98",X"C0",X"A9",X"00",X"85",X"73",X"20",
		X"44",X"B9",X"20",X"BA",X"C3",X"A9",X"A0",X"20",X"6A",X"B5",X"20",X"44",X"B9",X"A2",X"61",X"20",
		X"72",X"C7",X"20",X"55",X"B9",X"20",X"6C",X"DF",X"A5",X"37",X"29",X"07",X"C9",X"07",X"D0",X"02",
		X"A9",X"00",X"A8",X"84",X"9E",X"A9",X"08",X"20",X"4C",X"DF",X"A9",X"00",X"20",X"4A",X"DF",X"20",
		X"67",X"B9",X"20",X"39",X"DF",X"C6",X"37",X"10",X"AC",X"20",X"44",X"B9",X"A9",X"01",X"20",X"6A",
		X"DF",X"20",X"09",X"DF",X"A6",X"74",X"A4",X"75",X"A5",X"76",X"85",X"74",X"86",X"76",X"A5",X"77",
		X"85",X"75",X"84",X"77",X"60",X"A5",X"57",X"4A",X"4A",X"4A",X"4A",X"A0",X"00",X"C8",X"4A",X"D0",
		X"FC",X"18",X"69",X"02",X"A0",X"00",X"60",X"AD",X"15",X"04",X"F0",X"09",X"AD",X"6F",X"CE",X"AE",
		X"6E",X"CE",X"B8",X"50",X"06",X"AD",X"87",X"CE",X"AE",X"86",X"CE",X"60",X"F0",X"E7",X"CF",X"AA",
		X"80",X"56",X"31",X"19",X"10",X"19",X"31",X"56",X"80",X"AA",X"CF",X"E7",X"F0",X"F0",X"F0",X"B8",
		X"80",X"48",X"10",X"10",X"10",X"10",X"10",X"48",X"80",X"B8",X"F0",X"F0",X"F0",X"F0",X"B8",X"B8",
		X"80",X"48",X"48",X"10",X"10",X"10",X"48",X"48",X"80",X"B8",X"B8",X"F0",X"EC",X"D5",X"B1",X"90",
		X"70",X"4F",X"2B",X"14",X"14",X"2B",X"4F",X"70",X"90",X"B1",X"D5",X"EC",X"F0",X"C0",X"A0",X"94",
		X"6C",X"60",X"40",X"10",X"10",X"40",X"60",X"6C",X"94",X"A0",X"C0",X"F0",X"D9",X"C2",X"AC",X"97",
		X"80",X"69",X"52",X"3C",X"27",X"10",X"35",X"5A",X"80",X"A6",X"CA",X"F0",X"EA",X"E0",X"9C",X"80",
		X"64",X"20",X"16",X"50",X"16",X"20",X"64",X"80",X"9C",X"E0",X"EA",X"B0",X"10",X"1E",X"2C",X"3A",
		X"48",X"56",X"64",X"70",X"90",X"9E",X"AC",X"BA",X"C8",X"D6",X"E4",X"F0",X"10",X"1E",X"2D",X"3C",
		X"4B",X"5A",X"69",X"78",X"87",X"96",X"A5",X"B4",X"C3",X"D2",X"E1",X"F0",X"10",X"10",X"10",X"10",
		X"16",X"29",X"46",X"69",X"97",X"BA",X"D7",X"EA",X"F0",X"F0",X"F0",X"F0",X"10",X"24",X"30",X"36",
		X"3E",X"49",X"5A",X"75",X"94",X"A4",X"AC",X"BA",X"DA",X"E2",X"EA",X"F0",X"80",X"70",X"48",X"20",
		X"10",X"20",X"48",X"70",X"80",X"90",X"B8",X"E0",X"F0",X"E0",X"B8",X"90",X"DA",X"A4",X"87",X"80",
		X"79",X"5C",X"26",X"10",X"10",X"20",X"48",X"80",X"B8",X"E0",X"F0",X"F0",X"10",X"10",X"30",X"30",
		X"50",X"50",X"70",X"70",X"90",X"90",X"B0",X"B0",X"D0",X"D0",X"F0",X"F0",X"B0",X"80",X"50",X"47",
		X"18",X"30",X"18",X"47",X"50",X"80",X"B0",X"B9",X"E8",X"D4",X"E8",X"B9",X"10",X"1E",X"21",X"28",
		X"3C",X"55",X"66",X"73",X"8D",X"9A",X"AB",X"C4",X"D8",X"DF",X"E2",X"F0",X"80",X"AA",X"CF",X"E7",
		X"F0",X"E7",X"CF",X"AA",X"80",X"56",X"31",X"19",X"10",X"19",X"31",X"56",X"80",X"B8",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"B8",X"80",X"48",X"10",X"10",X"10",X"10",X"10",X"48",X"80",X"B8",X"B8",X"F0",
		X"F0",X"F0",X"B8",X"B8",X"80",X"48",X"48",X"10",X"10",X"10",X"48",X"48",X"94",X"B0",X"B8",X"A7",
		X"A7",X"B8",X"B0",X"94",X"6C",X"50",X"48",X"59",X"59",X"48",X"50",X"6C",X"96",X"A3",X"C5",X"F0",
		X"F0",X"C5",X"A3",X"96",X"6A",X"5D",X"3B",X"10",X"10",X"3B",X"5D",X"6A",X"3D",X"6A",X"97",X"C4",
		X"F0",X"C4",X"97",X"6A",X"3D",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"A0",X"E0",X"EA",X"B0",
		X"EA",X"E0",X"A0",X"80",X"60",X"20",X"16",X"50",X"16",X"20",X"60",X"80",X"F0",X"D0",X"B0",X"90",
		X"70",X"50",X"30",X"10",X"10",X"30",X"50",X"70",X"90",X"B0",X"D0",X"F0",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"F0",X"CB",X"A6",X"80",
		X"5C",X"39",X"20",X"12",X"12",X"20",X"39",X"5C",X"80",X"A6",X"CB",X"F0",X"C0",X"A6",X"8A",X"6A",
		X"4A",X"2F",X"14",X"24",X"20",X"39",X"59",X"75",X"72",X"90",X"B0",X"D0",X"80",X"57",X"48",X"57",
		X"80",X"A9",X"BA",X"A9",X"80",X"57",X"48",X"57",X"80",X"A9",X"BA",X"A9",X"E4",X"E8",X"B7",X"80",
		X"B7",X"E8",X"E4",X"B2",X"7A",X"47",X"20",X"10",X"20",X"47",X"7A",X"B2",X"90",X"70",X"70",X"50",
		X"50",X"30",X"30",X"10",X"10",X"30",X"30",X"50",X"50",X"70",X"70",X"90",X"E6",X"D0",X"E6",X"B9",
		X"AE",X"80",X"52",X"47",X"14",X"30",X"14",X"47",X"52",X"80",X"AE",X"B9",X"7E",X"6A",X"51",X"3A",
		X"2C",X"2C",X"38",X"4E",X"4E",X"38",X"2C",X"2C",X"3A",X"51",X"6A",X"7E",X"05",X"06",X"07",X"08",
		X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"00",X"01",X"02",X"03",X"04",X"04",X"04",X"08",X"08",
		X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"08",X"04",X"08",
		X"08",X"0C",X"08",X"0C",X"0C",X"00",X"0C",X"00",X"00",X"04",X"00",X"04",X"06",X"07",X"09",X"08",
		X"07",X"09",X"0A",X"0C",X"0E",X"0F",X"01",X"00",X"0F",X"01",X"02",X"04",X"07",X"06",X"05",X"08",
		X"0B",X"0A",X"09",X"0C",X"0F",X"0E",X"0D",X"00",X"03",X"02",X"01",X"04",X"05",X"05",X"05",X"05",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"04",X"08",X"0B",X"05",
		X"08",X"0C",X"0E",X"09",X"0C",X"00",X"03",X"0D",X"00",X"04",X"07",X"02",X"0D",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"0D",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0D",
		X"0E",X"0F",X"0F",X"00",X"01",X"01",X"02",X"03",X"04",X"04",X"04",X"00",X"0E",X"0D",X"0C",X"0D",
		X"0D",X"0D",X"01",X"0F",X"02",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"0B",X"09",X"07",X"05",
		X"03",X"01",X"0F",X"0D",X"0D",X"0F",X"01",X"03",X"05",X"07",X"09",X"0B",X"08",X"0B",X"0C",X"04",
		X"05",X"08",X"0B",X"0C",X"0D",X"0E",X"0F",X"01",X"02",X"03",X"04",X"05",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",X"0A",X"06",X"0C",X"08",
		X"0E",X"0A",X"00",X"0C",X"02",X"0E",X"04",X"00",X"06",X"02",X"08",X"04",X"0E",X"0C",X"0D",X"0E",
		X"00",X"02",X"02",X"00",X"0E",X"0E",X"00",X"02",X"03",X"04",X"02",X"00",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"0D",X"09",X"08",X"0C",X"0E",X"0F",X"0A",X"0B",X"18",X"1C",X"18",X"0F",
		X"18",X"18",X"18",X"18",X"0A",X"18",X"10",X"0F",X"18",X"0C",X"14",X"0A",X"50",X"50",X"50",X"68",
		X"50",X"50",X"68",X"B0",X"A0",X"50",X"90",X"80",X"20",X"B0",X"60",X"A0",X"40",X"20",X"40",X"80",
		X"40",X"40",X"70",X"60",X"00",X"20",X"40",X"00",X"A0",X"40",X"40",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"01",X"FF",X"00",X"00",X"FE",X"01",X"FF",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"60",X"40",
		X"00",X"00",X"48",X"40",X"50",X"28",X"50",X"00",X"00",X"50",X"00",X"40",X"04",X"04",X"03",X"04",
		X"04",X"04",X"03",X"04",X"05",X"04",X"04",X"04",X"04",X"04",X"04",X"05",X"3E",X"85",X"55",X"B9",
		X"35",X"04",X"85",X"56",X"B9",X"45",X"04",X"85",X"58",X"20",X"98",X"C0",X"A2",X"61",X"20",X"65",
		X"C7",X"A9",X"00",X"85",X"A9",X"20",X"3E",X"BD",X"A5",X"78",X"49",X"07",X"0A",X"C9",X"0A",X"B0",
		X"02",X"A9",X"0A",X"0A",X"0A",X"0A",X"0A",X"91",X"74",X"C8",X"A9",X"60",X"91",X"74",X"C8",X"84",
		X"A9",X"A4",X"55",X"BE",X"C9",X"CE",X"B9",X"C8",X"CE",X"A4",X"A9",X"4C",X"59",X"DF",X"A5",X"57",
		X"C9",X"10",X"90",X"48",X"38",X"E5",X"5F",X"8D",X"95",X"60",X"A9",X"00",X"E5",X"5B",X"8D",X"96",
		X"60",X"A9",X"18",X"8D",X"8C",X"60",X"A5",X"A0",X"8D",X"8E",X"60",X"8D",X"94",X"60",X"2C",X"40",
		X"60",X"30",X"FB",X"AD",X"60",X"60",X"85",X"79",X"AD",X"70",X"60",X"85",X"7A",X"A2",X"0F",X"8E",
		X"8C",X"60",X"38",X"E9",X"01",X"D0",X"02",X"A9",X"01",X"A2",X"00",X"E8",X"06",X"79",X"2A",X"90",
		X"FA",X"4A",X"49",X"7F",X"18",X"69",X"01",X"A8",X"8A",X"B8",X"50",X"04",X"A9",X"01",X"A0",X"00",
		X"85",X"78",X"48",X"98",X"A4",X"A9",X"91",X"74",X"C8",X"68",X"09",X"70",X"91",X"74",X"C8",X"60",
		X"85",X"36",X"B9",X"CE",X"03",X"85",X"56",X"B9",X"DE",X"03",X"85",X"58",X"A5",X"57",X"85",X"2F",
		X"98",X"18",X"69",X"01",X"29",X"0F",X"AA",X"BD",X"CE",X"03",X"85",X"2E",X"BD",X"DE",X"03",X"85",
		X"30",X"A9",X"00",X"85",X"59",X"A9",X"04",X"85",X"5A",X"A4",X"36",X"A5",X"5B",X"30",X"07",X"A5",
		X"57",X"C5",X"5F",X"B0",X"01",X"60",X"B9",X"B6",X"BF",X"85",X"99",X"B9",X"C4",X"BF",X"85",X"38",
		X"A4",X"9E",X"A9",X"08",X"20",X"4C",X"DF",X"20",X"98",X"C0",X"A2",X"61",X"20",X"65",X"C7",X"A5",
		X"2E",X"85",X"56",X"A5",X"2F",X"85",X"57",X"A5",X"30",X"85",X"58",X"20",X"98",X"C0",X"A4",X"59",
		X"A5",X"5A",X"20",X"6C",X"DF",X"A5",X"61",X"38",X"E5",X"6A",X"85",X"79",X"A5",X"62",X"E5",X"6B",
		X"85",X"9B",X"30",X"09",X"F0",X"04",X"A9",X"FF",X"85",X"79",X"B8",X"50",X"16",X"C9",X"FF",X"F0",
		X"05",X"A9",X"FF",X"B8",X"50",X"0B",X"A5",X"79",X"49",X"FF",X"18",X"69",X"01",X"90",X"02",X"A9",
		X"FF",X"85",X"79",X"A5",X"63",X"38",X"E5",X"6C",X"85",X"89",X"A5",X"64",X"E5",X"6D",X"85",X"9D",
		X"30",X"09",X"F0",X"04",X"A9",X"FF",X"85",X"89",X"B8",X"50",X"12",X"C9",X"FF",X"F0",X"05",X"A9",
		X"FF",X"B8",X"50",X"07",X"A5",X"89",X"49",X"FF",X"18",X"69",X"01",X"85",X"89",X"A9",X"00",X"85",
		X"82",X"85",X"92",X"A5",X"79",X"0A",X"26",X"82",X"85",X"7A",X"0A",X"85",X"7C",X"A5",X"82",X"2A",
		X"85",X"84",X"A5",X"7C",X"65",X"79",X"85",X"7D",X"A5",X"84",X"69",X"00",X"85",X"85",X"A5",X"7A",
		X"65",X"79",X"85",X"7B",X"A5",X"82",X"69",X"00",X"85",X"83",X"85",X"86",X"A5",X"7B",X"0A",X"85",
		X"7E",X"26",X"86",X"65",X"79",X"85",X"7F",X"A5",X"86",X"69",X"00",X"85",X"87",X"A5",X"89",X"0A",
		X"26",X"92",X"85",X"8A",X"0A",X"85",X"8C",X"A5",X"92",X"2A",X"85",X"94",X"A5",X"8C",X"65",X"89",
		X"85",X"8D",X"A5",X"94",X"69",X"00",X"85",X"95",X"A5",X"8A",X"65",X"89",X"85",X"8B",X"A5",X"92",
		X"69",X"00",X"85",X"93",X"85",X"96",X"A5",X"8B",X"0A",X"85",X"8E",X"26",X"96",X"65",X"89",X"85",
		X"8F",X"A5",X"96",X"69",X"00",X"85",X"97",X"A0",X"00",X"84",X"A9",X"A4",X"38",X"B9",X"D3",X"BF",
		X"C9",X"01",X"D0",X"02",X"A9",X"C0",X"85",X"73",X"B9",X"D2",X"BF",X"85",X"2D",X"C8",X"C8",X"84",
		X"38",X"AA",X"29",X"07",X"A8",X"8A",X"0A",X"85",X"2B",X"4A",X"4A",X"4A",X"4A",X"29",X"07",X"AA",
		X"A5",X"2B",X"45",X"9B",X"30",X"0B",X"B9",X"78",X"00",X"85",X"61",X"B9",X"80",X"00",X"B8",X"50",
		X"11",X"B9",X"78",X"00",X"49",X"FF",X"18",X"69",X"01",X"85",X"61",X"B9",X"80",X"00",X"49",X"FF",
		X"69",X"00",X"85",X"62",X"A5",X"2D",X"45",X"9D",X"10",X"0E",X"B5",X"88",X"18",X"65",X"61",X"85",
		X"61",X"B5",X"90",X"65",X"62",X"B8",X"50",X"0B",X"A5",X"61",X"38",X"F5",X"88",X"85",X"61",X"A5",
		X"62",X"F5",X"90",X"85",X"62",X"A5",X"2B",X"45",X"9D",X"30",X"0B",X"B9",X"88",X"00",X"85",X"63",
		X"B9",X"90",X"00",X"B8",X"50",X"11",X"B9",X"88",X"00",X"49",X"FF",X"18",X"69",X"01",X"85",X"63",
		X"B9",X"90",X"00",X"49",X"FF",X"69",X"00",X"85",X"64",X"A5",X"2D",X"45",X"9B",X"10",X"0E",X"A5",
		X"63",X"38",X"F5",X"78",X"85",X"63",X"A5",X"64",X"F5",X"80",X"B8",X"50",X"0B",X"A5",X"63",X"18",
		X"75",X"78",X"85",X"63",X"A5",X"64",X"75",X"80",X"85",X"64",X"A4",X"A9",X"A5",X"63",X"91",X"74",
		X"C8",X"A5",X"64",X"29",X"1F",X"91",X"74",X"C8",X"A5",X"61",X"91",X"74",X"C8",X"A5",X"62",X"29",
		X"1F",X"05",X"73",X"91",X"74",X"C8",X"84",X"A9",X"C6",X"99",X"F0",X"03",X"4C",X"DB",X"BE",X"A4",
		X"A9",X"88",X"4C",X"5F",X"DF",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"06",
		X"07",X"07",X"04",X"02",X"00",X"10",X"20",X"30",X"40",X"50",X"60",X"70",X"80",X"92",X"9E",X"AC",
		X"BA",X"C2",X"0C",X"01",X"8C",X"01",X"4A",X"01",X"09",X"01",X"CB",X"01",X"4B",X"01",X"89",X"01",
		X"CA",X"01",X"90",X"01",X"8A",X"01",X"23",X"01",X"DB",X"01",X"41",X"01",X"10",X"01",X"0A",X"01",
		X"CB",X"01",X"91",X"01",X"17",X"01",X"4B",X"01",X"8A",X"01",X"CE",X"01",X"08",X"01",X"0A",X"01",
		X"CB",X"01",X"92",X"01",X"16",X"01",X"4B",X"01",X"8A",X"01",X"CD",X"01",X"49",X"01",X"0A",X"01",
		X"CB",X"01",X"93",X"01",X"15",X"01",X"4B",X"01",X"8A",X"01",X"CC",X"01",X"4A",X"01",X"0A",X"01",
		X"CB",X"01",X"95",X"01",X"13",X"01",X"4B",X"01",X"8A",X"01",X"CA",X"01",X"4C",X"01",X"0A",X"01",
		X"CB",X"01",X"96",X"01",X"12",X"01",X"4B",X"01",X"8A",X"01",X"C9",X"01",X"4D",X"01",X"0A",X"01",
		X"CB",X"01",X"97",X"01",X"11",X"01",X"4B",X"01",X"8A",X"01",X"88",X"01",X"4E",X"01",X"0A",X"01",
		X"CB",X"01",X"0B",X"00",X"A3",X"01",X"0A",X"01",X"10",X"01",X"4B",X"01",X"8A",X"01",X"90",X"01",
		X"41",X"01",X"5B",X"01",X"9A",X"01",X"31",X"01",X"B1",X"01",X"31",X"01",X"B1",X"01",X"1A",X"01",
		X"01",X"00",X"91",X"01",X"21",X"01",X"A1",X"01",X"21",X"01",X"A1",X"01",X"11",X"01",X"01",X"00",
		X"89",X"01",X"11",X"01",X"91",X"01",X"11",X"01",X"91",X"01",X"09",X"01",X"01",X"00",X"8A",X"01",
		X"12",X"01",X"8A",X"01",X"01",X"00",X"06",X"01",X"A5",X"57",X"38",X"E5",X"5F",X"8D",X"95",X"60",
		X"A9",X"00",X"E5",X"5B",X"8D",X"96",X"60",X"10",X"0A",X"A9",X"00",X"8D",X"96",X"60",X"A9",X"01",
		X"8D",X"95",X"60",X"A5",X"58",X"C5",X"60",X"90",X"07",X"E5",X"60",X"A2",X"00",X"B8",X"50",X"07",
		X"A5",X"60",X"38",X"E5",X"58",X"A2",X"FF",X"8D",X"8E",X"60",X"8D",X"94",X"60",X"86",X"33",X"A5",
		X"56",X"C5",X"5E",X"90",X"07",X"E5",X"5E",X"A2",X"00",X"B8",X"50",X"07",X"A5",X"5E",X"38",X"E5",
		X"56",X"A2",X"FF",X"85",X"32",X"86",X"34",X"2C",X"40",X"60",X"30",X"FB",X"AD",X"60",X"60",X"85",
		X"63",X"AD",X"70",X"60",X"85",X"64",X"A5",X"32",X"8D",X"8E",X"60",X"8D",X"94",X"60",X"A5",X"33",
		X"30",X"18",X"A5",X"63",X"18",X"65",X"68",X"85",X"63",X"A5",X"64",X"65",X"69",X"50",X"06",X"A9",
		X"FF",X"85",X"63",X"A9",X"7F",X"85",X"64",X"B8",X"50",X"15",X"A5",X"68",X"38",X"E5",X"63",X"85",
		X"63",X"A5",X"69",X"E5",X"64",X"50",X"06",X"A9",X"00",X"85",X"63",X"A9",X"80",X"85",X"64",X"2C",
		X"40",X"60",X"30",X"FB",X"AD",X"60",X"60",X"85",X"61",X"AD",X"70",X"60",X"85",X"62",X"A6",X"34",
		X"30",X"16",X"A5",X"61",X"18",X"65",X"66",X"85",X"61",X"A5",X"62",X"65",X"67",X"50",X"06",X"A9",
		X"FF",X"85",X"61",X"A9",X"7F",X"85",X"62",X"60",X"A5",X"66",X"38",X"E5",X"61",X"85",X"61",X"A5",
		X"67",X"E5",X"62",X"50",X"06",X"A9",X"00",X"85",X"61",X"A9",X"80",X"85",X"62",X"60",X"20",X"13",
		X"AA",X"A9",X"80",X"85",X"5E",X"A9",X"FF",X"8D",X"14",X"01",X"20",X"35",X"C2",X"AD",X"33",X"01",
		X"D0",X"03",X"8D",X"00",X"58",X"A9",X"00",X"8D",X"33",X"01",X"AD",X"C6",X"CE",X"8D",X"00",X"20",
		X"AD",X"C7",X"CE",X"8D",X"01",X"20",X"A5",X"9F",X"29",X"70",X"C9",X"5F",X"90",X"02",X"A9",X"5F",
		X"4A",X"09",X"07",X"AA",X"A0",X"07",X"BD",X"FD",X"C1",X"29",X"0F",X"99",X"19",X"00",X"99",X"00",
		X"08",X"BD",X"FD",X"C1",X"4A",X"4A",X"4A",X"4A",X"99",X"21",X"00",X"99",X"08",X"08",X"CA",X"88",
		X"10",X"E4",X"60",X"A9",X"00",X"85",X"81",X"85",X"91",X"85",X"80",X"85",X"78",X"85",X"90",X"85",
		X"88",X"A9",X"00",X"8D",X"80",X"60",X"8D",X"81",X"60",X"8D",X"84",X"60",X"8D",X"85",X"60",X"8D",
		X"86",X"60",X"8D",X"87",X"60",X"8D",X"89",X"60",X"8D",X"83",X"60",X"8D",X"8D",X"60",X"8D",X"8E",
		X"60",X"8D",X"8F",X"60",X"8D",X"90",X"60",X"A9",X"0F",X"8D",X"8C",X"60",X"60",X"00",X"04",X"08",
		X"0C",X"C3",X"07",X"0B",X"0B",X"00",X"07",X"0B",X"08",X"44",X"03",X"0C",X"0C",X"00",X"0B",X"03",
		X"07",X"C8",X"0C",X"04",X"04",X"00",X"0B",X"08",X"07",X"C4",X"0C",X"03",X"03",X"00",X"04",X"08",
		X"0C",X"C3",X"07",X"0F",X"0B",X"00",X"0C",X"08",X"04",X"C3",X"0B",X"07",X"07",X"06",X"03",X"01",
		X"04",X"00",X"05",X"05",X"05",X"A6",X"3D",X"B5",X"46",X"20",X"E8",X"C2",X"48",X"AC",X"12",X"01",
		X"B9",X"8C",X"BC",X"49",X"FF",X"18",X"69",X"01",X"85",X"5F",X"85",X"5D",X"A9",X"10",X"38",X"E5",
		X"5F",X"85",X"A0",X"A9",X"FF",X"85",X"5B",X"B9",X"9C",X"BC",X"85",X"60",X"B9",X"CC",X"BC",X"8D",
		X"11",X"01",X"A5",X"02",X"C9",X"1E",X"D0",X"0D",X"B9",X"AC",X"BC",X"85",X"68",X"B9",X"BC",X"BC",
		X"85",X"69",X"B8",X"50",X"18",X"B9",X"AC",X"BC",X"38",X"E5",X"68",X"8D",X"21",X"01",X"B9",X"BC",
		X"BC",X"ED",X"69",X"00",X"A2",X"03",X"4A",X"6E",X"21",X"01",X"CA",X"10",X"F9",X"A9",X"00",X"85",
		X"66",X"85",X"67",X"A9",X"00",X"8D",X"0F",X"01",X"8D",X"10",X"01",X"A9",X"2C",X"8D",X"13",X"01",
		X"68",X"A8",X"A2",X"0F",X"B9",X"7C",X"B9",X"9D",X"CE",X"03",X"B9",X"7C",X"BA",X"9D",X"DE",X"03",
		X"A9",X"00",X"9D",X"1A",X"03",X"9D",X"3A",X"03",X"9D",X"9A",X"03",X"B9",X"7C",X"BB",X"9D",X"EE",
		X"03",X"88",X"CA",X"10",X"DF",X"A0",X"00",X"A2",X"0F",X"B9",X"CE",X"03",X"38",X"7D",X"CE",X"03",
		X"6A",X"9D",X"35",X"04",X"B9",X"DE",X"03",X"38",X"7D",X"DE",X"03",X"6A",X"9D",X"45",X"04",X"88",
		X"10",X"02",X"A0",X"0F",X"CA",X"10",X"E2",X"60",X"A2",X"00",X"C9",X"62",X"90",X"05",X"AD",X"CA",
		X"60",X"29",X"5F",X"C9",X"10",X"90",X"04",X"E8",X"38",X"E9",X"10",X"C9",X"10",X"B0",X"F6",X"A8",
		X"B9",X"7C",X"BC",X"8D",X"12",X"01",X"0A",X"0A",X"0A",X"0A",X"09",X"0F",X"60",X"AD",X"10",X"01",
		X"D0",X"27",X"A9",X"F0",X"85",X"57",X"A2",X"4F",X"20",X"73",X"C4",X"8D",X"10",X"01",X"F0",X"03",
		X"8D",X"0F",X"01",X"AD",X"0F",X"01",X"D0",X"11",X"A9",X"10",X"85",X"57",X"20",X"53",X"C4",X"A5",
		X"57",X"A2",X"0F",X"20",X"73",X"C4",X"8D",X"0F",X"01",X"A9",X"01",X"20",X"6A",X"DF",X"A0",X"06",
		X"84",X"9E",X"AE",X"10",X"01",X"F0",X"01",X"60",X"AE",X"13",X"01",X"D0",X"01",X"60",X"A2",X"0F",
		X"A9",X"C0",X"20",X"EE",X"C3",X"CA",X"10",X"F8",X"A0",X"06",X"84",X"9E",X"A9",X"08",X"20",X"4C",
		X"DF",X"A0",X"4F",X"AD",X"10",X"01",X"20",X"6E",X"C3",X"A0",X"0F",X"AD",X"0F",X"01",X"D0",X"49",
		X"84",X"37",X"B9",X"2A",X"03",X"85",X"61",X"B9",X"1A",X"03",X"85",X"62",X"B9",X"4A",X"03",X"85",
		X"63",X"B9",X"3A",X"03",X"85",X"64",X"A2",X"61",X"20",X"72",X"C7",X"A5",X"74",X"85",X"B0",X"A5",
		X"75",X"85",X"B1",X"A2",X"0F",X"AD",X"11",X"01",X"F0",X"01",X"CA",X"A9",X"C0",X"85",X"73",X"86",
		X"38",X"C6",X"37",X"A5",X"37",X"29",X"0F",X"C9",X"0F",X"D0",X"07",X"A5",X"37",X"18",X"69",X"10",
		X"85",X"37",X"20",X"23",X"C4",X"C6",X"38",X"10",X"E8",X"60",X"A5",X"61",X"38",X"E5",X"6A",X"85",
		X"6E",X"A5",X"62",X"E5",X"6B",X"85",X"6F",X"A5",X"63",X"38",X"E5",X"6C",X"85",X"70",X"A5",X"64",
		X"E5",X"6D",X"85",X"71",X"A2",X"6E",X"20",X"92",X"DF",X"A5",X"61",X"85",X"6A",X"A5",X"62",X"85",
		X"6B",X"A5",X"63",X"85",X"6C",X"A5",X"64",X"85",X"6D",X"A9",X"C0",X"85",X"73",X"60",X"86",X"37",
		X"48",X"A4",X"9E",X"A9",X"08",X"20",X"4C",X"DF",X"20",X"3C",X"C4",X"A2",X"61",X"20",X"72",X"C7",
		X"68",X"85",X"73",X"48",X"20",X"23",X"C4",X"C6",X"37",X"A4",X"9E",X"A9",X"00",X"85",X"73",X"A9",
		X"08",X"20",X"4C",X"DF",X"20",X"23",X"C4",X"68",X"85",X"73",X"20",X"3C",X"C4",X"20",X"BA",X"C3",
		X"A6",X"37",X"60",X"A6",X"37",X"BD",X"2A",X"03",X"85",X"61",X"BD",X"1A",X"03",X"85",X"62",X"BD",
		X"4A",X"03",X"85",X"63",X"BD",X"3A",X"03",X"85",X"64",X"4C",X"BA",X"C3",X"A6",X"37",X"BD",X"6A",
		X"03",X"85",X"61",X"BD",X"5A",X"03",X"85",X"62",X"BD",X"8A",X"03",X"85",X"63",X"BD",X"7A",X"03",
		X"85",X"64",X"60",X"A5",X"5B",X"D0",X"1A",X"A5",X"57",X"38",X"E5",X"5F",X"90",X"02",X"C9",X"0C",
		X"B0",X"0F",X"A5",X"5F",X"18",X"69",X"0F",X"B0",X"02",X"C9",X"F0",X"90",X"02",X"A9",X"F0",X"85",
		X"57",X"60",X"DB",X"85",X"57",X"86",X"38",X"A9",X"00",X"85",X"59",X"A2",X"0F",X"86",X"37",X"A6",
		X"37",X"BD",X"CE",X"03",X"85",X"56",X"BD",X"DE",X"03",X"85",X"58",X"20",X"98",X"C0",X"A6",X"38",
		X"A4",X"61",X"A5",X"62",X"30",X"0D",X"C9",X"04",X"90",X"06",X"A0",X"FF",X"A9",X"03",X"E6",X"59",
		X"B8",X"50",X"0A",X"C9",X"FC",X"B0",X"06",X"A0",X"01",X"A9",X"FC",X"E6",X"59",X"9D",X"1A",X"03",
		X"98",X"9D",X"2A",X"03",X"A4",X"63",X"A5",X"64",X"30",X"0D",X"C9",X"04",X"90",X"06",X"A0",X"FF",
		X"A9",X"03",X"E6",X"59",X"B8",X"50",X"0A",X"C9",X"FC",X"B0",X"06",X"A9",X"FC",X"A0",X"01",X"E6",
		X"59",X"9D",X"3A",X"03",X"98",X"9D",X"4A",X"03",X"C6",X"38",X"C6",X"37",X"10",X"A1",X"A5",X"59",
		X"60",X"20",X"E8",X"C2",X"85",X"36",X"86",X"35",X"A9",X"00",X"85",X"73",X"A9",X"05",X"20",X"6A",
		X"DF",X"A5",X"35",X"29",X"07",X"AA",X"BC",X"2D",X"C2",X"84",X"9E",X"A9",X"08",X"20",X"4C",X"DF",
		X"AE",X"12",X"01",X"A5",X"36",X"BC",X"CC",X"BC",X"D0",X"03",X"38",X"E9",X"0F",X"A8",X"B9",X"7C",
		X"BA",X"85",X"57",X"49",X"80",X"AA",X"B9",X"7C",X"B9",X"85",X"56",X"49",X"80",X"20",X"75",X"DF",
		X"A9",X"C0",X"85",X"73",X"A2",X"0F",X"86",X"38",X"A4",X"36",X"B9",X"7C",X"B9",X"AA",X"38",X"E5",
		X"56",X"48",X"86",X"56",X"B9",X"7C",X"BA",X"A8",X"38",X"E5",X"57",X"AA",X"84",X"57",X"68",X"20",
		X"75",X"DF",X"C6",X"36",X"C6",X"38",X"10",X"E0",X"A9",X"01",X"4C",X"6A",X"DF",X"AD",X"15",X"01",
		X"F0",X"5F",X"A5",X"5F",X"48",X"A5",X"5B",X"48",X"A5",X"A0",X"48",X"A9",X"E8",X"85",X"5F",X"A9",
		X"FF",X"85",X"5B",X"A9",X"28",X"85",X"A0",X"A2",X"07",X"86",X"37",X"A6",X"37",X"BD",X"FE",X"03",
		X"F0",X"32",X"85",X"57",X"A9",X"80",X"85",X"56",X"A9",X"80",X"85",X"58",X"A5",X"9F",X"C9",X"05",
		X"B0",X"05",X"A9",X"06",X"B8",X"50",X"09",X"8A",X"29",X"07",X"C9",X"07",X"D0",X"02",X"A9",X"04",
		X"85",X"9E",X"A8",X"A9",X"08",X"20",X"4C",X"DF",X"A5",X"37",X"29",X"03",X"0A",X"69",X"0A",X"85",
		X"55",X"20",X"09",X"BD",X"C6",X"37",X"10",X"C3",X"68",X"85",X"A0",X"68",X"85",X"5B",X"68",X"85",
		X"5F",X"AD",X"1F",X"01",X"F0",X"0B",X"A6",X"42",X"E0",X"15",X"90",X"05",X"A6",X"40",X"FE",X"00",
		X"02",X"60",X"AD",X"10",X"01",X"F0",X"01",X"60",X"A5",X"5B",X"D0",X"07",X"A5",X"5F",X"C9",X"F0",
		X"90",X"01",X"60",X"A9",X"01",X"20",X"6A",X"DF",X"A5",X"74",X"48",X"A5",X"75",X"48",X"A9",X"00",
		X"85",X"38",X"85",X"A9",X"A2",X"0F",X"AD",X"11",X"01",X"F0",X"01",X"CA",X"86",X"37",X"A2",X"03",
		X"A4",X"A9",X"BD",X"69",X"C6",X"91",X"74",X"C8",X"CA",X"10",X"F7",X"84",X"A9",X"AD",X"14",X"01",
		X"D0",X"4A",X"A6",X"38",X"BD",X"9A",X"03",X"30",X"11",X"A2",X"0B",X"A4",X"A9",X"B1",X"AA",X"91",
		X"74",X"C8",X"CA",X"10",X"F8",X"84",X"A9",X"B8",X"50",X"2F",X"A4",X"A9",X"B1",X"AA",X"91",X"74",
		X"85",X"6C",X"C8",X"B1",X"AA",X"91",X"74",X"C9",X"10",X"90",X"02",X"09",X"E0",X"85",X"6D",X"C8",
		X"B1",X"AA",X"91",X"74",X"85",X"6A",X"C8",X"B1",X"AA",X"91",X"74",X"C9",X"10",X"90",X"02",X"09",
		X"E0",X"85",X"6B",X"C8",X"84",X"A9",X"20",X"C7",X"C6",X"B8",X"50",X"06",X"20",X"6D",X"C6",X"20",
		X"C7",X"C6",X"A6",X"38",X"1E",X"9A",X"03",X"E6",X"38",X"C6",X"37",X"10",X"91",X"68",X"85",X"AB",
		X"68",X"85",X"AA",X"A4",X"A9",X"88",X"4C",X"5F",X"DF",X"80",X"40",X"68",X"05",X"A5",X"38",X"AA",
		X"18",X"69",X"01",X"29",X"0F",X"A8",X"BD",X"6A",X"03",X"38",X"79",X"6A",X"03",X"85",X"61",X"BD",
		X"5A",X"03",X"79",X"5A",X"03",X"85",X"62",X"0A",X"66",X"62",X"66",X"61",X"BD",X"8A",X"03",X"38",
		X"79",X"8A",X"03",X"85",X"63",X"BD",X"7A",X"03",X"79",X"7A",X"03",X"85",X"64",X"0A",X"66",X"64",
		X"66",X"63",X"A4",X"A9",X"A5",X"63",X"91",X"74",X"C8",X"85",X"6C",X"A5",X"64",X"85",X"6D",X"29",
		X"1F",X"91",X"74",X"C8",X"A5",X"61",X"91",X"74",X"C8",X"85",X"6A",X"A5",X"62",X"85",X"6B",X"29",
		X"1F",X"91",X"74",X"C8",X"84",X"A9",X"60",X"A6",X"38",X"BD",X"AC",X"03",X"D0",X"16",X"A4",X"A9",
		X"A2",X"03",X"A9",X"00",X"91",X"74",X"C8",X"A9",X"71",X"91",X"74",X"C8",X"CA",X"10",X"F3",X"84",
		X"A9",X"B8",X"50",X"57",X"85",X"57",X"20",X"53",X"C4",X"BD",X"35",X"04",X"85",X"56",X"BD",X"45",
		X"04",X"85",X"58",X"20",X"98",X"C0",X"20",X"3C",X"C7",X"A6",X"38",X"BD",X"9A",X"03",X"29",X"40",
		X"F0",X"1F",X"20",X"3E",X"BD",X"AD",X"CA",X"60",X"29",X"02",X"18",X"69",X"1C",X"AA",X"BD",X"C9",
		X"CE",X"C8",X"91",X"74",X"88",X"BD",X"C8",X"CE",X"91",X"74",X"C8",X"C8",X"84",X"A9",X"B8",X"50",
		X"1A",X"A4",X"A9",X"A9",X"00",X"91",X"74",X"C8",X"A9",X"68",X"91",X"74",X"C8",X"AD",X"B2",X"3D",
		X"91",X"74",X"C8",X"AD",X"B3",X"3D",X"91",X"74",X"C8",X"84",X"A9",X"60",X"A4",X"A9",X"A5",X"63",
		X"38",X"E5",X"6C",X"91",X"74",X"C8",X"A5",X"64",X"E5",X"6D",X"29",X"1F",X"91",X"74",X"C8",X"A5",
		X"61",X"38",X"E5",X"6A",X"91",X"74",X"C8",X"A5",X"62",X"E5",X"6B",X"29",X"1F",X"09",X"A0",X"91",
		X"74",X"C8",X"84",X"A9",X"60",X"A0",X"00",X"98",X"91",X"74",X"A9",X"71",X"C8",X"91",X"74",X"C8",
		X"D0",X"02",X"A0",X"00",X"A9",X"40",X"91",X"74",X"A9",X"80",X"C8",X"91",X"74",X"C8",X"B5",X"02",
		X"85",X"6C",X"91",X"74",X"C8",X"B5",X"03",X"85",X"6D",X"29",X"1F",X"91",X"74",X"B5",X"00",X"85",
		X"6A",X"C8",X"91",X"74",X"B5",X"01",X"85",X"6B",X"29",X"1F",X"C8",X"91",X"74",X"4C",X"5F",X"DF",
		X"20",X"95",X"CD",X"A9",X"00",X"85",X"00",X"A5",X"53",X"C9",X"09",X"90",X"FA",X"A9",X"00",X"85",
		X"53",X"20",X"BD",X"C7",X"20",X"91",X"C8",X"20",X"B6",X"B1",X"18",X"90",X"EA",X"AD",X"00",X"0D",
		X"29",X"83",X"C9",X"82",X"F0",X"13",X"20",X"D2",X"A7",X"A6",X"00",X"A5",X"4E",X"09",X"80",X"85",
		X"4E",X"BD",X"DB",X"C7",X"48",X"BD",X"DA",X"C7",X"48",X"60",X"0B",X"C9",X"3F",X"C9",X"0A",X"97",
		X"AE",X"C9",X"F0",X"C9",X"FF",X"C7",X"00",X"00",X"8B",X"C9",X"3E",X"AC",X"6D",X"AD",X"17",X"CA",
		X"48",X"91",X"4A",X"90",X"E6",X"B0",X"07",X"91",X"7A",X"C9",X"28",X"97",X"E0",X"D7",X"17",X"A6",
		X"E6",X"06",X"85",X"17",X"A5",X"07",X"4A",X"B0",X"27",X"A0",X"00",X"A2",X"02",X"B5",X"13",X"F0",
		X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",X"95",X"13",X"CA",X"10",X"F0",X"98",X"D0",X"10",
		X"A2",X"02",X"B5",X"13",X"F0",X"07",X"18",X"69",X"EF",X"95",X"13",X"30",X"03",X"CA",X"10",X"F2",
		X"60",X"5D",X"D1",X"8F",X"D1",X"8F",X"D1",X"B1",X"D1",X"EB",X"D1",X"03",X"D2",X"61",X"D2",X"CB",
		X"D2",X"33",X"D3",X"66",X"D3",X"B0",X"D3",X"E6",X"D3",X"FF",X"D3",X"17",X"D4",X"1D",X"D4",X"34",
		X"D4",X"4C",X"D4",X"60",X"D4",X"A1",X"D4",X"AB",X"D4",X"EF",X"D4",X"30",X"D5",X"75",X"D5",X"85",
		X"D5",X"A1",X"D5",X"A8",X"D5",X"E9",X"D5",X"1C",X"D6",X"62",X"D6",X"7A",X"D6",X"67",X"D1",X"97",
		X"D1",X"97",X"D1",X"BD",X"D1",X"F0",X"D1",X"17",X"D2",X"75",X"D2",X"E0",X"D2",X"3F",X"D3",X"79",
		X"D3",X"BE",X"D3",X"E6",X"D3",X"FF",X"D3",X"17",X"D4",X"22",X"D4",X"3A",X"D4",X"51",X"D4",X"6D",
		X"D4",X"A1",X"D4",X"BA",X"D4",X"FD",X"D4",X"3F",X"D5",X"75",X"D5",X"85",X"D5",X"A1",X"D5",X"B9",
		X"D5",X"F6",X"D5",X"29",X"D6",X"68",X"D6",X"7A",X"D6",X"75",X"D1",X"9F",X"D1",X"9F",X"D1",X"CF",
		X"D1",X"F6",X"D1",X"30",X"D2",X"94",X"D2",X"FB",X"D2",X"50",X"D3",X"8B",X"D3",X"CB",X"D3",X"F5",
		X"D3",X"0E",X"D4",X"17",X"D4",X"28",X"D4",X"41",X"D4",X"5B",X"D4",X"83",X"D4",X"A1",X"D4",X"CC",
		X"D4",X"0E",X"D5",X"51",X"D5",X"75",X"D5",X"8E",X"D5",X"A1",X"D5",X"C8",X"D5",X"04",X"D6",X"3E",
		X"D6",X"6F",X"D6",X"8F",X"D6",X"7F",X"D1",X"A8",X"D1",X"A8",X"D1",X"DE",X"D1",X"FC",X"D1",X"4D",
		X"D2",X"AE",X"D2",X"16",X"D3",X"5E",X"D3",X"A0",X"D3",X"DA",X"D3",X"ED",X"D3",X"06",X"D4",X"17",
		X"D4",X"2D",X"D4",X"46",X"D4",X"56",X"D4",X"92",X"D4",X"A1",X"D4",X"DD",X"D4",X"1F",X"D5",X"63",
		X"D5",X"75",X"D5",X"97",X"D5",X"A1",X"D5",X"D9",X"D5",X"10",X"D6",X"51",X"D6",X"74",X"D6",X"A1",
		X"D6",X"51",X"56",X"00",X"1A",X"01",X"20",X"31",X"56",X"01",X"38",X"31",X"B0",X"41",X"00",X"11",
		X"F6",X"30",X"38",X"31",X"CE",X"51",X"0A",X"31",X"E2",X"31",X"E2",X"51",X"BA",X"51",X"98",X"51",
		X"D8",X"51",X"C9",X"31",X"56",X"51",X"80",X"51",X"80",X"51",X"80",X"51",X"80",X"71",X"92",X"51",
		X"80",X"31",X"B0",X"51",X"89",X"41",X"89",X"00",X"00",X"71",X"5A",X"71",X"A0",X"E5",X"22",X"16",
		X"2E",X"1E",X"00",X"32",X"40",X"1E",X"B8",X"D9",X"20",X"26",X"30",X"00",X"1C",X"1E",X"00",X"34",
		X"16",X"38",X"3C",X"26",X"9E",X"E5",X"3A",X"34",X"26",X"1E",X"2C",X"1E",X"30",X"1C",X"9E",X"D3",
		X"28",X"3E",X"1E",X"22",X"32",X"00",X"3C",X"1E",X"38",X"2E",X"26",X"30",X"16",X"1C",X"B2",X"CD",
		X"34",X"2C",X"16",X"46",X"1E",X"38",X"80",X"C6",X"28",X"32",X"3E",X"1E",X"3E",X"38",X"80",X"C6",
		X"3A",X"34",X"26",X"1E",X"2C",X"1E",X"38",X"80",X"C6",X"28",X"3E",X"22",X"16",X"1C",X"32",X"38",
		X"80",X"DF",X"34",X"38",X"1E",X"3A",X"3A",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"CD",X"16",X"34",
		X"34",X"3E",X"46",X"1E",X"48",X"00",X"3A",X"3E",X"38",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"D6",
		X"3A",X"3C",X"16",X"38",X"3C",X"00",X"1C",X"38",X"3E",X"1E",X"1A",X"2A",X"1E",X"B0",X"DC",X"34",
		X"3E",X"2C",X"3A",X"16",X"38",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"F4",X"34",X"2C",X"16",X"C6",
		X"F1",X"28",X"32",X"3E",X"1E",X"C8",X"F1",X"3A",X"34",X"26",X"1E",X"AC",X"EE",X"28",X"3E",X"1E",
		X"22",X"3E",X"9E",X"C7",X"1E",X"30",X"3C",X"1E",X"38",X"00",X"46",X"32",X"3E",X"38",X"00",X"26",
		X"30",X"26",X"3C",X"26",X"16",X"2C",X"BA",X"B8",X"3A",X"40",X"34",X"00",X"1E",X"30",X"3C",X"38",
		X"1E",X"48",X"00",X"40",X"32",X"3A",X"00",X"26",X"30",X"26",X"3C",X"26",X"16",X"2C",X"1E",X"BA",
		X"AC",X"22",X"1E",X"18",X"1E",X"30",X"00",X"3A",X"26",X"1E",X"00",X"26",X"24",X"38",X"1E",X"00",
		X"26",X"30",X"26",X"3C",X"26",X"16",X"2C",X"1E",X"30",X"00",X"1E",X"26",X"B0",X"C7",X"1E",X"30",
		X"3C",X"38",X"1E",X"00",X"3A",X"3E",X"3A",X"00",X"26",X"30",X"26",X"1A",X"26",X"16",X"2C",X"1E",
		X"BA",X"C7",X"3A",X"34",X"26",X"30",X"00",X"2A",X"30",X"32",X"18",X"00",X"3C",X"32",X"00",X"1A",
		X"24",X"16",X"30",X"22",X"9E",X"A6",X"3C",X"32",X"3E",X"38",X"30",X"1E",X"48",X"00",X"2C",X"1E",
		X"00",X"18",X"32",X"3E",X"3C",X"32",X"30",X"00",X"34",X"32",X"3E",X"38",X"00",X"1A",X"24",X"16",
		X"30",X"22",X"1E",X"B8",X"B5",X"2A",X"30",X"32",X"34",X"20",X"00",X"1C",X"38",X"1E",X"24",X"1E",
		X"30",X"00",X"48",X"3E",X"2E",X"00",X"42",X"1E",X"1A",X"24",X"3A",X"1E",X"2C",X"B0",X"AC",X"22",
		X"26",X"38",X"1E",X"00",X"2C",X"16",X"00",X"34",X"1E",X"38",X"26",X"2C",X"2C",X"16",X"00",X"34",
		X"16",X"38",X"16",X"00",X"1A",X"16",X"2E",X"18",X"26",X"16",X"B8",X"C4",X"34",X"38",X"1E",X"3A",
		X"3A",X"00",X"20",X"26",X"38",X"1E",X"00",X"3C",X"32",X"00",X"3A",X"1E",X"2C",X"1E",X"1A",X"BC",
		X"B2",X"34",X"32",X"3E",X"3A",X"3A",X"1E",X"48",X"00",X"20",X"1E",X"3E",X"00",X"36",X"3E",X"16",
		X"30",X"1C",X"00",X"1A",X"32",X"38",X"38",X"1E",X"1A",X"3C",X"9E",X"B2",X"20",X"26",X"38",X"1E",
		X"00",X"1C",X"38",X"3E",X"1E",X"1A",X"2A",X"1E",X"30",X"00",X"42",X"1E",X"30",X"30",X"00",X"38",
		X"26",X"1A",X"24",X"3C",X"26",X"A2",X"AC",X"32",X"34",X"38",X"26",X"2E",X"16",X"00",X"20",X"26",
		X"38",X"1E",X"00",X"34",X"16",X"38",X"16",X"00",X"3A",X"1E",X"2C",X"1E",X"1A",X"1A",X"26",X"32",
		X"30",X"16",X"B8",X"BC",X"24",X"26",X"22",X"24",X"00",X"3A",X"1A",X"32",X"38",X"1E",X"BA",X"9E",
		X"2E",X"1E",X"26",X"2C",X"2C",X"1E",X"3E",X"38",X"3A",X"00",X"3A",X"1A",X"32",X"38",X"1E",X"BA",
		X"B0",X"24",X"32",X"1E",X"1A",X"24",X"3A",X"3C",X"48",X"16",X"24",X"2C",X"1E",X"B0",X"D4",X"38",
		X"1E",X"1A",X"32",X"38",X"1C",X"BA",X"C2",X"38",X"16",X"30",X"2A",X"26",X"30",X"22",X"00",X"20",
		X"38",X"32",X"2E",X"00",X"04",X"00",X"3C",X"32",X"80",X"C2",X"34",X"2C",X"16",X"1A",X"1E",X"2E",
		X"1E",X"30",X"3C",X"00",X"1C",X"1E",X"00",X"04",X"00",X"16",X"80",X"BC",X"38",X"16",X"30",X"22",
		X"2C",X"26",X"3A",X"3C",X"1E",X"00",X"40",X"32",X"30",X"00",X"04",X"00",X"48",X"3E",X"2E",X"80",
		X"C8",X"38",X"16",X"30",X"2A",X"26",X"30",X"22",X"00",X"1C",X"1E",X"00",X"04",X"00",X"16",X"80",
		X"D9",X"38",X"16",X"3C",X"1E",X"00",X"46",X"32",X"3E",X"38",X"3A",X"1E",X"2C",X"A0",X"DC",X"1E",
		X"40",X"16",X"2C",X"3E",X"1E",X"48",X"4C",X"40",X"32",X"3E",X"BA",X"D6",X"3A",X"1E",X"2C",X"18",
		X"3A",X"3C",X"00",X"38",X"1E",X"1A",X"24",X"30",X"1E",X"B0",X"DF",X"1A",X"16",X"2C",X"26",X"20",
		X"26",X"36",X"3E",X"1E",X"3A",X"9E",X"AA",X"30",X"32",X"40",X"26",X"1A",X"9E",X"AA",X"30",X"32",
		X"40",X"26",X"1A",X"26",X"B2",X"AA",X"16",X"30",X"20",X"16",X"1E",X"30",X"22",X"1E",X"B8",X"4A",
		X"1E",X"44",X"34",X"1E",X"38",X"BC",X"45",X"1E",X"44",X"34",X"1E",X"38",X"3C",X"B2",X"40",X"1E",
		X"38",X"20",X"16",X"24",X"38",X"1E",X"B0",X"8B",X"18",X"32",X"30",X"3E",X"BA",X"E8",X"3C",X"26",
		X"2E",X"9E",X"E0",X"1C",X"3E",X"38",X"1E",X"9E",X"E8",X"48",X"1E",X"26",X"BC",X"E4",X"3C",X"26",
		X"1E",X"2E",X"34",X"B2",X"8B",X"2C",X"1E",X"40",X"1E",X"AC",X"8B",X"30",X"26",X"40",X"1E",X"16",
		X"BE",X"8B",X"22",X"38",X"16",X"9C",X"8B",X"30",X"26",X"40",X"1E",X"AC",X"8B",X"24",X"32",X"2C",
		X"9E",X"8B",X"3C",X"38",X"32",X"BE",X"8B",X"24",X"32",X"46",X"B2",X"8B",X"2C",X"32",X"1A",X"A4",
		X"DC",X"26",X"30",X"3A",X"1E",X"38",X"3C",X"00",X"1A",X"32",X"26",X"30",X"BA",X"C1",X"26",X"30",
		X"3C",X"38",X"32",X"1C",X"3E",X"26",X"38",X"1E",X"00",X"2C",X"1E",X"3A",X"00",X"34",X"26",X"1E",
		X"1A",X"1E",X"BA",X"D6",X"22",X"1E",X"2C",X"1C",X"00",X"1E",X"26",X"30",X"42",X"1E",X"38",X"20",
		X"1E",X"B0",X"D6",X"26",X"30",X"3A",X"1E",X"38",X"3C",X"1E",X"00",X"20",X"26",X"1A",X"24",X"16",
		X"BA",X"00",X"20",X"38",X"1E",X"1E",X"00",X"34",X"2C",X"16",X"C6",X"0E",X"04",X"00",X"1A",X"32",
		X"26",X"30",X"00",X"06",X"00",X"34",X"2C",X"16",X"46",X"BA",X"FA",X"04",X"00",X"34",X"26",X"1E",
		X"1A",X"1E",X"00",X"06",X"00",X"28",X"32",X"3E",X"1E",X"3E",X"38",X"BA",X"00",X"04",X"00",X"2E",
		X"3E",X"1E",X"30",X"48",X"00",X"06",X"00",X"3A",X"34",X"26",X"1E",X"2C",X"9E",X"FA",X"04",X"00",
		X"2E",X"32",X"30",X"1E",X"1C",X"16",X"00",X"06",X"00",X"28",X"3E",X"1E",X"22",X"32",X"BA",X"14",
		X"04",X"00",X"1A",X"32",X"26",X"30",X"00",X"04",X"00",X"34",X"2C",X"16",X"C6",X"00",X"04",X"00",
		X"34",X"26",X"1E",X"1A",X"1E",X"00",X"04",X"00",X"28",X"32",X"3E",X"1E",X"3E",X"B8",X"00",X"04",
		X"00",X"2E",X"3E",X"1E",X"30",X"48",X"1E",X"00",X"04",X"00",X"3A",X"34",X"26",X"1E",X"AC",X"00",
		X"04",X"00",X"2E",X"32",X"30",X"1E",X"1C",X"16",X"00",X"04",X"00",X"28",X"3E",X"1E",X"22",X"B2",
		X"0E",X"06",X"00",X"1A",X"32",X"26",X"30",X"3A",X"00",X"04",X"00",X"34",X"2C",X"16",X"C6",X"FA",
		X"06",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"3A",X"00",X"04",X"00",X"28",X"32",X"3E",X"1E",X"3E",
		X"B8",X"FA",X"06",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"1E",X"30",X"00",X"04",X"00",X"3A",X"34",
		X"26",X"1E",X"AC",X"FA",X"06",X"00",X"2E",X"32",X"30",X"1E",X"1C",X"16",X"3A",X"00",X"04",X"00",
		X"28",X"3E",X"1E",X"22",X"B2",X"D3",X"50",X"00",X"2E",X"1A",X"2E",X"2C",X"44",X"44",X"44",X"00",
		X"16",X"3C",X"16",X"38",X"A6",X"A0",X"1A",X"38",X"1E",X"1C",X"26",X"3C",X"3A",X"80",X"A0",X"2A",
		X"38",X"1E",X"1C",X"26",X"3C",X"1E",X"80",X"A0",X"1A",X"38",X"1E",X"1C",X"26",X"3C",X"32",X"3A",
		X"80",X"DA",X"18",X"32",X"30",X"3E",X"3A",X"80",X"D0",X"06",X"00",X"1A",X"38",X"1E",X"1C",X"26",
		X"3C",X"00",X"2E",X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D6",X"06",X"00",X"28",X"1E",X"3E",X"44",
		X"00",X"2E",X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D0",X"06",X"00",X"3A",X"34",X"26",X"1E",X"2C",
		X"1E",X"00",X"2E",X"26",X"30",X"26",X"2E",X"3E",X"AE",X"D3",X"06",X"00",X"28",X"3E",X"1E",X"22",
		X"32",X"3A",X"00",X"2E",X"26",X"30",X"26",X"2E",X"B2",X"C8",X"18",X"32",X"30",X"3E",X"3A",X"00",
		X"1E",X"40",X"1E",X"38",X"46",X"80",X"CE",X"18",X"32",X"30",X"3E",X"3A",X"00",X"1A",X"24",X"16",
		X"36",X"3E",X"1E",X"80",X"CE",X"18",X"32",X"30",X"3E",X"3A",X"00",X"28",X"1E",X"1C",X"1E",X"80",
		X"C8",X"18",X"32",X"30",X"3E",X"3A",X"00",X"1A",X"16",X"1C",X"16",X"80",X"B8",X"16",X"40",X"32",
		X"26",X"1C",X"00",X"3A",X"34",X"26",X"2A",X"1E",X"BA",X"88",X"16",X"3C",X"3C",X"1E",X"30",X"3C",
		X"26",X"32",X"30",X"00",X"16",X"3E",X"44",X"00",X"2C",X"16",X"30",X"1A",X"1E",X"BA",X"96",X"3A",
		X"34",X"26",X"3C",X"48",X"1E",X"30",X"00",X"16",X"3E",X"3A",X"42",X"1E",X"26",X"1A",X"24",X"1E",
		X"B0",X"A0",X"1E",X"40",X"26",X"3C",X"1E",X"00",X"2C",X"16",X"3A",X"00",X"34",X"3E",X"30",X"3C",
		X"16",X"BA",X"E0",X"2C",X"1E",X"40",X"1E",X"AC",X"DA",X"30",X"26",X"40",X"1E",X"16",X"BE",X"E2",
		X"22",X"38",X"16",X"9C",X"E0",X"30",X"26",X"40",X"1E",X"AC",X"C4",X"3A",X"3E",X"34",X"1E",X"38",
		X"48",X"16",X"34",X"34",X"1E",X"38",X"00",X"38",X"1E",X"1A",X"24",X"16",X"38",X"22",X"9E",X"CD",
		X"30",X"1E",X"3E",X"1E",X"38",X"00",X"3A",X"3E",X"34",X"1E",X"38",X"48",X"16",X"34",X"34",X"1E",
		X"B8",X"CD",X"30",X"3E",X"1E",X"40",X"32",X"00",X"3A",X"3E",X"34",X"1E",X"38",X"48",X"16",X"34",
		X"34",X"1E",X"B8",X"31",X"D0",X"6D",X"D0",X"A9",X"D0",X"E5",X"D0",X"AD",X"00",X"0E",X"85",X"0A",
		X"29",X"38",X"4A",X"4A",X"4A",X"AA",X"BD",X"F7",X"D6",X"8D",X"56",X"01",X"AD",X"00",X"0D",X"49",
		X"02",X"85",X"09",X"A5",X"0A",X"2A",X"2A",X"2A",X"29",X"03",X"AA",X"BD",X"FF",X"D6",X"8D",X"58",
		X"01",X"A5",X"0A",X"29",X"06",X"A8",X"B9",X"B3",X"D6",X"85",X"AC",X"B9",X"B4",X"D6",X"85",X"AD",
		X"20",X"E0",X"DB",X"8D",X"6A",X"01",X"60",X"02",X"01",X"03",X"04",X"05",X"06",X"07",X"00",X"03",
		X"04",X"05",X"02",X"7C",X"48",X"8A",X"48",X"98",X"48",X"D8",X"BA",X"E0",X"D0",X"90",X"04",X"A5",
		X"53",X"10",X"04",X"00",X"4C",X"3F",X"D9",X"8D",X"00",X"50",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"49",X"0F",X"A8",X"29",X"10",X"8D",X"17",X"01",X"98",X"38",X"E5",X"52",X"29",X"0F",X"C9",X"08",
		X"90",X"02",X"09",X"F0",X"18",X"65",X"50",X"85",X"50",X"84",X"52",X"8D",X"DB",X"60",X"AC",X"D8",
		X"60",X"AD",X"00",X"0C",X"85",X"08",X"A5",X"4C",X"84",X"4C",X"A8",X"25",X"4C",X"05",X"4D",X"85",
		X"4D",X"98",X"05",X"4C",X"25",X"4D",X"85",X"4D",X"A8",X"45",X"4F",X"25",X"4D",X"05",X"4E",X"85",
		X"4E",X"84",X"4F",X"A5",X"B4",X"A4",X"13",X"10",X"02",X"09",X"04",X"A4",X"14",X"10",X"02",X"09",
		X"02",X"A4",X"15",X"10",X"02",X"09",X"01",X"8D",X"00",X"40",X"A6",X"3E",X"E8",X"A4",X"05",X"D0",
		X"10",X"A2",X"00",X"A4",X"07",X"C0",X"40",X"90",X"08",X"A6",X"06",X"E0",X"02",X"90",X"02",X"A2",
		X"03",X"BD",X"DD",X"D7",X"45",X"A1",X"29",X"03",X"45",X"A1",X"85",X"A1",X"8D",X"E0",X"60",X"20",
		X"24",X"CF",X"20",X"0A",X"CD",X"E6",X"53",X"E6",X"07",X"D0",X"1E",X"EE",X"06",X"04",X"D0",X"08",
		X"EE",X"07",X"04",X"D0",X"03",X"EE",X"08",X"04",X"24",X"05",X"50",X"0D",X"EE",X"09",X"04",X"D0",
		X"08",X"EE",X"0A",X"04",X"D0",X"03",X"EE",X"0B",X"04",X"2C",X"00",X"0C",X"50",X"09",X"EE",X"33",
		X"01",X"8D",X"00",X"58",X"8D",X"00",X"48",X"68",X"A8",X"68",X"AA",X"68",X"40",X"FF",X"FD",X"FE",
		X"FC",X"A9",X"00",X"85",X"05",X"A9",X"02",X"85",X"01",X"AD",X"CA",X"01",X"D0",X"15",X"AD",X"00",
		X"0C",X"29",X"10",X"F0",X"0E",X"A9",X"00",X"85",X"00",X"AD",X"C9",X"01",X"29",X"03",X"F0",X"03",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7",
		X"20",X"AC",X"AB",X"60",X"20",X"BB",X"D6",X"20",X"A8",X"AA",X"20",X"0D",X"DD",X"20",X"41",X"DD",
		X"AD",X"58",X"01",X"85",X"37",X"20",X"53",X"DF",X"A9",X"E8",X"A2",X"C0",X"20",X"75",X"DF",X"A9",
		X"32",X"A2",X"6C",X"20",X"39",X"DF",X"C6",X"37",X"D0",X"F5",X"AD",X"6A",X"01",X"29",X"03",X"0A",
		X"A8",X"B9",X"1F",X"3F",X"BE",X"1E",X"3F",X"20",X"39",X"DF",X"AD",X"00",X"02",X"20",X"CE",X"AD",
		X"8D",X"00",X"02",X"29",X"06",X"48",X"A8",X"B9",X"17",X"3F",X"BE",X"16",X"3F",X"20",X"39",X"DF",
		X"68",X"4A",X"AA",X"A5",X"4D",X"3D",X"B6",X"D8",X"DD",X"B6",X"D8",X"D0",X"1A",X"CA",X"CA",X"10",
		X"03",X"4C",X"3F",X"D9",X"D0",X"06",X"20",X"E9",X"DD",X"B8",X"50",X"0B",X"20",X"ED",X"DD",X"AD",
		X"C9",X"01",X"09",X"03",X"8D",X"C9",X"01",X"AD",X"CA",X"01",X"2D",X"C6",X"01",X"F0",X"07",X"A9",
		X"34",X"A2",X"6E",X"20",X"39",X"DF",X"20",X"53",X"DF",X"A5",X"09",X"29",X"1C",X"4A",X"4A",X"AA",
		X"BD",X"BA",X"D8",X"A0",X"EE",X"A2",X"1B",X"20",X"A9",X"D8",X"A5",X"09",X"4A",X"4A",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"C2",X"D8",X"A0",X"32",X"A2",X"F8",X"85",X"29",X"98",X"20",X"75",X"DF",X"A9",
		X"29",X"A0",X"01",X"4C",X"B1",X"DF",X"18",X"18",X"30",X"50",X"11",X"14",X"15",X"16",X"21",X"24",
		X"25",X"26",X"00",X"12",X"14",X"24",X"15",X"13",X"00",X"00",X"A8",X"A9",X"00",X"84",X"79",X"4A",
		X"4A",X"0A",X"AA",X"98",X"29",X"0F",X"D0",X"01",X"E8",X"9A",X"A9",X"A2",X"8D",X"C1",X"60",X"BA",
		X"D0",X"07",X"A9",X"60",X"A0",X"09",X"B8",X"50",X"04",X"A9",X"C0",X"A0",X"01",X"8D",X"C0",X"60",
		X"A9",X"03",X"8D",X"E0",X"60",X"A2",X"00",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",
		X"FB",X"8D",X"00",X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",X"C1",X"60",X"A9",X"00",X"8D",
		X"E0",X"60",X"A0",X"09",X"2C",X"00",X"0C",X"30",X"FB",X"2C",X"00",X"0C",X"10",X"FB",X"8D",X"00",
		X"50",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"BA",X"CA",X"9A",X"10",X"AE",X"4C",X"0A",X"DA",X"51",
		X"00",X"A8",X"A5",X"01",X"C9",X"20",X"90",X"02",X"E9",X"18",X"29",X"1F",X"4C",X"CD",X"D8",X"78",
		X"8D",X"00",X"50",X"8D",X"00",X"58",X"A2",X"FF",X"9A",X"D8",X"E8",X"8A",X"A8",X"84",X"00",X"86",
		X"01",X"A0",X"00",X"91",X"00",X"C8",X"D0",X"FB",X"E8",X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",
		X"30",X"8D",X"00",X"50",X"90",X"E7",X"85",X"01",X"8D",X"E0",X"60",X"8D",X"CF",X"60",X"8D",X"DF",
		X"60",X"A2",X"07",X"8E",X"CF",X"60",X"8E",X"DF",X"60",X"E8",X"9D",X"C0",X"60",X"9D",X"D0",X"60",
		X"CA",X"10",X"F7",X"AD",X"00",X"0C",X"29",X"10",X"F0",X"1F",X"8D",X"00",X"50",X"CE",X"00",X"01",
		X"D0",X"F8",X"CE",X"01",X"01",X"D0",X"F3",X"A9",X"10",X"85",X"B4",X"20",X"11",X"DE",X"20",X"AC",
		X"AB",X"20",X"6E",X"C1",X"58",X"4C",X"A0",X"C7",X"A0",X"A2",X"11",X"9A",X"A0",X"00",X"BA",X"96",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"F0",X"03",X"4C",X"CA",X"D8",X"E8",X"D0",X"F4",X"BA",
		X"8A",X"8D",X"00",X"50",X"C8",X"59",X"00",X"00",X"D0",X"EF",X"99",X"00",X"00",X"C8",X"D0",X"DE",
		X"BA",X"8A",X"0A",X"AA",X"90",X"D5",X"A0",X"00",X"A2",X"01",X"84",X"00",X"86",X"01",X"A0",X"00",
		X"B1",X"00",X"F0",X"03",X"4C",X"31",X"D9",X"A9",X"11",X"91",X"00",X"D1",X"00",X"F0",X"03",X"4C",
		X"2F",X"D9",X"0A",X"90",X"F4",X"A9",X"00",X"91",X"00",X"C8",X"D0",X"E4",X"8D",X"00",X"50",X"E8",
		X"E0",X"08",X"D0",X"02",X"A2",X"20",X"E0",X"30",X"90",X"D0",X"A9",X"00",X"A8",X"AA",X"85",X"3B",
		X"A9",X"30",X"85",X"3C",X"A9",X"08",X"85",X"38",X"8A",X"51",X"3B",X"C8",X"D0",X"FB",X"E6",X"3C",
		X"8D",X"00",X"50",X"C6",X"38",X"D0",X"F2",X"95",X"7D",X"E8",X"E0",X"02",X"D0",X"04",X"A9",X"90",
		X"85",X"3C",X"E0",X"0C",X"90",X"DE",X"A5",X"7D",X"F0",X"0A",X"A9",X"40",X"A2",X"A4",X"8D",X"C4",
		X"60",X"8E",X"C5",X"60",X"A2",X"05",X"AD",X"CA",X"60",X"CD",X"CA",X"60",X"D0",X"05",X"CA",X"10",
		X"F8",X"85",X"7A",X"A2",X"05",X"AD",X"DA",X"60",X"CD",X"DA",X"60",X"D0",X"05",X"CA",X"10",X"F8",
		X"85",X"7B",X"20",X"11",X"DE",X"A0",X"02",X"AD",X"C9",X"01",X"F0",X"0A",X"85",X"7C",X"20",X"F1",
		X"DD",X"A0",X"00",X"8C",X"C9",X"01",X"84",X"00",X"A2",X"07",X"BD",X"F9",X"DA",X"9D",X"00",X"08",
		X"CA",X"10",X"F7",X"A9",X"00",X"8D",X"E0",X"60",X"A9",X"10",X"8D",X"00",X"40",X"A0",X"04",X"A2",
		X"14",X"2C",X"00",X"0C",X"10",X"FB",X"2C",X"00",X"0C",X"30",X"FB",X"CA",X"10",X"F3",X"88",X"30",
		X"08",X"8D",X"00",X"50",X"2C",X"00",X"0C",X"50",X"E6",X"8D",X"00",X"58",X"A9",X"00",X"85",X"74",
		X"A9",X"20",X"85",X"75",X"8D",X"CB",X"60",X"AD",X"C8",X"60",X"85",X"52",X"29",X"0F",X"85",X"50",
		X"AD",X"00",X"0C",X"49",X"FF",X"29",X"2F",X"85",X"4E",X"29",X"28",X"F0",X"0B",X"06",X"4C",X"90",
		X"04",X"E6",X"00",X"E6",X"00",X"B8",X"50",X"04",X"A9",X"20",X"85",X"4C",X"20",X"0F",X"DB",X"20",
		X"0D",X"DF",X"8D",X"00",X"48",X"E6",X"03",X"A5",X"03",X"29",X"03",X"D0",X"03",X"20",X"1B",X"DE",
		X"AD",X"00",X"0C",X"29",X"10",X"F0",X"96",X"D0",X"FE",X"00",X"04",X"08",X"0C",X"03",X"07",X"0B",
		X"0B",X"59",X"DB",X"F6",X"DB",X"83",X"DB",X"99",X"DB",X"7D",X"DB",X"6E",X"DB",X"21",X"DB",X"A6",
		X"00",X"E0",X"0E",X"90",X"04",X"A2",X"02",X"86",X"00",X"BD",X"02",X"DB",X"48",X"BD",X"01",X"DB",
		X"48",X"60",X"A9",X"00",X"8D",X"E0",X"60",X"8D",X"80",X"60",X"8D",X"C0",X"60",X"8D",X"D0",X"60",
		X"8D",X"00",X"60",X"8D",X"40",X"60",X"AD",X"40",X"60",X"AD",X"60",X"60",X"AD",X"70",X"60",X"AD",
		X"50",X"60",X"A9",X"08",X"8D",X"E0",X"60",X"A9",X"01",X"A2",X"1F",X"18",X"9D",X"80",X"60",X"2A",
		X"CA",X"10",X"F9",X"A9",X"34",X"A2",X"A6",X"4C",X"39",X"DF",X"AD",X"CA",X"01",X"0D",X"C7",X"01",
		X"D0",X"0C",X"20",X"11",X"DE",X"AD",X"C9",X"01",X"85",X"7C",X"A9",X"02",X"85",X"00",X"60",X"A5",
		X"50",X"4A",X"A8",X"A9",X"68",X"20",X"4C",X"DF",X"A2",X"4E",X"A9",X"33",X"D0",X"0A",X"A2",X"B6",
		X"A9",X"32",X"D0",X"04",X"A9",X"33",X"A2",X"0A",X"20",X"39",X"DF",X"A2",X"06",X"A9",X"00",X"9D",
		X"C1",X"60",X"9D",X"D1",X"60",X"CA",X"CA",X"10",X"F6",X"60",X"A5",X"03",X"29",X"3F",X"D0",X"02",
		X"E6",X"39",X"A5",X"39",X"29",X"07",X"AA",X"BC",X"D5",X"DB",X"A9",X"00",X"99",X"C1",X"60",X"BC",
		X"D6",X"DB",X"BD",X"DC",X"DF",X"99",X"C0",X"60",X"A9",X"A8",X"99",X"C1",X"60",X"A9",X"34",X"A2",
		X"56",X"20",X"39",X"DF",X"A5",X"03",X"29",X"7F",X"A8",X"A9",X"01",X"20",X"6C",X"DF",X"A9",X"34",
		X"A2",X"AA",X"4C",X"39",X"DF",X"16",X"00",X"10",X"02",X"12",X"04",X"14",X"06",X"16",X"00",X"EA",
		X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"07",X"85",X"37",X"8D",X"CB",X"60",X"AD",X"C8",X"60",
		X"29",X"20",X"4A",X"4A",X"05",X"37",X"60",X"A5",X"2E",X"F0",X"1E",X"8D",X"95",X"60",X"8D",X"8D",
		X"60",X"A5",X"2F",X"8D",X"96",X"60",X"A2",X"00",X"20",X"E6",X"DC",X"C9",X"01",X"D0",X"06",X"98",
		X"D0",X"03",X"8A",X"10",X"04",X"A9",X"FF",X"85",X"78",X"A2",X"00",X"86",X"73",X"E6",X"2E",X"D0",
		X"06",X"E6",X"2F",X"10",X"02",X"86",X"2F",X"8D",X"DB",X"60",X"AD",X"D8",X"60",X"29",X"78",X"85",
		X"4D",X"F0",X"05",X"8D",X"C0",X"60",X"A2",X"A4",X"8E",X"C1",X"60",X"A2",X"00",X"A5",X"4E",X"F0",
		X"06",X"0A",X"8D",X"C2",X"60",X"A2",X"A4",X"8E",X"C3",X"60",X"20",X"0D",X"DD",X"A4",X"4D",X"A9",
		X"D0",X"A2",X"F0",X"20",X"2B",X"DD",X"A4",X"4E",X"20",X"27",X"DD",X"A5",X"52",X"29",X"10",X"F0",
		X"1D",X"A9",X"34",X"A2",X"82",X"20",X"39",X"DF",X"A0",X"10",X"A5",X"4D",X"29",X"60",X"F0",X"0E",
		X"49",X"20",X"F0",X"04",X"A9",X"04",X"A0",X"08",X"8D",X"E0",X"60",X"8C",X"00",X"40",X"A9",X"34",
		X"A2",X"92",X"20",X"39",X"DF",X"A2",X"0B",X"B5",X"7D",X"F0",X"19",X"85",X"35",X"86",X"38",X"8A",
		X"20",X"1F",X"DF",X"A0",X"F4",X"A2",X"F4",X"A5",X"35",X"20",X"A9",X"D8",X"A9",X"0C",X"AA",X"20",
		X"75",X"DF",X"A6",X"38",X"CA",X"10",X"E0",X"20",X"53",X"DF",X"A9",X"00",X"A2",X"16",X"20",X"75",
		X"DF",X"A2",X"04",X"86",X"37",X"A6",X"37",X"A0",X"00",X"B5",X"78",X"F0",X"03",X"BC",X"E1",X"DC",
		X"B9",X"E4",X"31",X"BE",X"E5",X"31",X"20",X"57",X"DF",X"C6",X"37",X"10",X"E8",X"A2",X"AC",X"A9",
		X"30",X"20",X"75",X"DF",X"A4",X"50",X"B9",X"E8",X"DF",X"BE",X"E4",X"DF",X"A0",X"C0",X"4C",X"73",
		X"DF",X"2E",X"38",X"34",X"36",X"1E",X"A0",X"00",X"84",X"73",X"8C",X"14",X"04",X"8D",X"8E",X"60",
		X"8E",X"8F",X"60",X"8C",X"90",X"60",X"A2",X"10",X"8E",X"8C",X"60",X"8E",X"94",X"60",X"CA",X"30",
		X"0B",X"AD",X"40",X"60",X"30",X"F8",X"AD",X"60",X"60",X"AC",X"70",X"60",X"60",X"20",X"53",X"DF",
		X"A9",X"00",X"20",X"6A",X"DF",X"A9",X"E8",X"AC",X"00",X"0D",X"20",X"29",X"DD",X"AC",X"00",X"0E",
		X"20",X"27",X"DD",X"20",X"E0",X"DB",X"A8",X"A9",X"D0",X"A2",X"F8",X"84",X"35",X"20",X"75",X"DF",
		X"A2",X"07",X"86",X"37",X"06",X"35",X"A9",X"00",X"2A",X"20",X"1F",X"DF",X"C6",X"37",X"10",X"F4",
		X"60",X"AD",X"0F",X"04",X"0A",X"85",X"29",X"AD",X"10",X"04",X"2A",X"85",X"2A",X"AD",X"0C",X"04",
		X"18",X"65",X"29",X"8D",X"95",X"60",X"85",X"29",X"AD",X"0D",X"04",X"65",X"2A",X"8D",X"96",X"60",
		X"05",X"29",X"D0",X"05",X"A9",X"01",X"8D",X"95",X"60",X"AD",X"09",X"04",X"8D",X"8D",X"60",X"AD",
		X"0A",X"04",X"AE",X"0B",X"04",X"20",X"E6",X"DC",X"8D",X"12",X"04",X"8C",X"13",X"04",X"A9",X"3D",
		X"A2",X"CE",X"20",X"39",X"DF",X"A9",X"06",X"85",X"3B",X"A9",X"04",X"85",X"3C",X"85",X"37",X"A0",
		X"00",X"84",X"31",X"84",X"32",X"84",X"33",X"84",X"34",X"B1",X"3B",X"85",X"56",X"E6",X"3B",X"B1",
		X"3B",X"85",X"57",X"E6",X"3B",X"B1",X"3B",X"85",X"58",X"E6",X"3B",X"F8",X"A0",X"17",X"84",X"38",
		X"26",X"56",X"26",X"57",X"26",X"58",X"A0",X"03",X"A2",X"00",X"B5",X"31",X"75",X"31",X"95",X"31",
		X"E8",X"88",X"10",X"F6",X"C6",X"38",X"10",X"E8",X"D8",X"A9",X"31",X"A0",X"04",X"20",X"B1",X"DF",
		X"A9",X"D0",X"A2",X"F8",X"20",X"75",X"DF",X"C6",X"37",X"10",X"B4",X"60",X"73",X"00",X"09",X"0A",
		X"15",X"16",X"22",X"15",X"06",X"15",X"07",X"06",X"04",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",
		X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",X"03",X"D0",X"02",X"A9",X"04",X"A0",X"00",X"8C",
		X"C6",X"01",X"48",X"0D",X"C7",X"01",X"8D",X"C7",X"01",X"68",X"0D",X"C8",X"01",X"8D",X"C8",X"01",
		X"60",X"A9",X"07",X"8D",X"C7",X"01",X"A9",X"00",X"8D",X"C8",X"01",X"AD",X"CA",X"01",X"D0",X"4B",
		X"AD",X"C7",X"01",X"F0",X"46",X"A2",X"00",X"8E",X"CB",X"01",X"8E",X"CF",X"01",X"8E",X"CE",X"01",
		X"A2",X"08",X"38",X"6E",X"CE",X"01",X"0A",X"CA",X"90",X"F9",X"A0",X"80",X"AD",X"CE",X"01",X"2D",
		X"C8",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"CA",X"01",X"AD",X"CE",X"01",X"4D",X"C7",X"01",X"8D",
		X"C7",X"01",X"8A",X"0A",X"AA",X"BD",X"DD",X"DD",X"8D",X"CC",X"01",X"BD",X"DE",X"DD",X"8D",X"CD",
		X"01",X"BD",X"E3",X"DD",X"85",X"BD",X"BD",X"E4",X"DD",X"85",X"BE",X"A0",X"00",X"8C",X"40",X"60",
		X"AD",X"CA",X"01",X"D0",X"01",X"60",X"AC",X"CB",X"01",X"AE",X"CC",X"01",X"0A",X"90",X"0D",X"9D",
		X"00",X"60",X"A9",X"40",X"8D",X"CA",X"01",X"A0",X"0E",X"B8",X"50",X"73",X"10",X"25",X"A9",X"80",
		X"8D",X"CA",X"01",X"AD",X"C6",X"01",X"F0",X"04",X"A9",X"00",X"91",X"BD",X"B1",X"BD",X"EC",X"CD",
		X"01",X"90",X"08",X"A9",X"00",X"8D",X"CA",X"01",X"AD",X"CF",X"01",X"9D",X"00",X"60",X"A0",X"0C",
		X"B8",X"50",X"3F",X"A9",X"08",X"8D",X"40",X"60",X"9D",X"00",X"60",X"A9",X"09",X"8D",X"40",X"60",
		X"EA",X"A9",X"08",X"8D",X"40",X"60",X"EC",X"CD",X"01",X"AD",X"50",X"60",X"90",X"20",X"4D",X"CF",
		X"01",X"F0",X"13",X"A9",X"00",X"AC",X"CB",X"01",X"91",X"BD",X"88",X"10",X"FB",X"AD",X"CE",X"01",
		X"0D",X"C9",X"01",X"8D",X"C9",X"01",X"A9",X"00",X"8D",X"CA",X"01",X"B8",X"50",X"02",X"91",X"BD",
		X"A0",X"00",X"18",X"6D",X"CF",X"01",X"8D",X"CF",X"01",X"EE",X"CB",X"01",X"EE",X"CC",X"01",X"8C",
		X"40",X"60",X"98",X"D0",X"03",X"4C",X"1B",X"DE",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"53",X"DF",
		X"A9",X"20",X"A0",X"00",X"91",X"74",X"4C",X"AC",X"DF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"E4",X"31",X"91",X"74",X"BD",X"E5",
		X"31",X"C8",X"91",X"74",X"20",X"5F",X"DF",X"28",X"60",X"4A",X"29",X"0F",X"09",X"A0",X"A0",X"01",
		X"91",X"74",X"88",X"8A",X"6A",X"91",X"74",X"C8",X"D0",X"15",X"A4",X"73",X"09",X"60",X"AA",X"98",
		X"4C",X"57",X"DF",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",X"74",X"C8",X"8A",X"91",X"74",X"98",
		X"38",X"65",X"74",X"85",X"74",X"90",X"02",X"E6",X"75",X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",
		X"4C",X"57",X"DF",X"84",X"73",X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"6F",X"0A",X"26",X"6F",
		X"85",X"6E",X"8A",X"0A",X"A0",X"00",X"90",X"01",X"88",X"84",X"71",X"0A",X"26",X"71",X"85",X"70",
		X"A2",X"6E",X"A0",X"00",X"B5",X"02",X"91",X"74",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"74",X"B5",
		X"00",X"C8",X"91",X"74",X"B5",X"01",X"45",X"73",X"29",X"1F",X"45",X"73",X"C8",X"91",X"74",X"D0",
		X"AE",X"38",X"08",X"88",X"84",X"AE",X"18",X"65",X"AE",X"28",X"AA",X"08",X"86",X"AF",X"B5",X"00",
		X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"19",X"DF",X"A5",X"AE",X"D0",X"01",X"18",X"A6",X"AF",X"B5",
		X"00",X"20",X"19",X"DF",X"A6",X"AF",X"CA",X"C6",X"AE",X"10",X"E0",X"60",X"10",X"10",X"40",X"40",
		X"90",X"90",X"FF",X"FF",X"00",X"0C",X"16",X"1E",X"20",X"1E",X"16",X"0C",X"00",X"F4",X"EA",X"E2",
		X"E0",X"E2",X"EA",X"F4",X"00",X"0C",X"16",X"1E",X"00",X"00",X"04",X"D7",X"3F",X"D9",X"04",X"D7");
begin
process(clk)
begin
	if rising_edge(clk) then
       if (clk_en) then
			data <= rom_data(to_integer(unsigned(addr)));
			end if;
	end if;
end process;
end architecture;
