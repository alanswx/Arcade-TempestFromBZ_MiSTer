module progrom
(
input clk,
input [14:0] addr,
output [7:0] dout,
input cs );
reg [7:0] q;
always @(posedge clk) 
begin 
case (addr) 
	15'h0: q<=8'h02;
	15'h1: q<=8'hbb;
	15'h2: q<=8'h5a;
	15'h3: q<=8'h30;
	15'h4: q<=8'h50;
	15'h5: q<=8'hee;
	15'h6: q<=8'h3d;
	15'h7: q<=8'ha8;
	15'h8: q<=8'h4d;
	15'h9: q<=8'h20;
	15'ha: q<=8'hc5;
	15'hb: q<=8'h92;
	15'hc: q<=8'h20;
	15'hd: q<=8'h34;
	15'he: q<=8'h92;
	15'hf: q<=8'h20;
	15'h10: q<=8'h2b;
	15'h11: q<=8'h90;
	15'h12: q<=8'h20;
	15'h13: q<=8'h31;
	15'h14: q<=8'ha8;
	15'h15: q<=8'ha9;
	15'h16: q<=8'hfa;
	15'h17: q<=8'h85;
	15'h18: q<=8'h5b;
	15'h19: q<=8'ha9;
	15'h1a: q<=8'h00;
	15'h1b: q<=8'h8d;
	15'h1c: q<=8'h06;
	15'h1d: q<=8'h01;
	15'h1e: q<=8'h85;
	15'h1f: q<=8'h5f;
	15'h20: q<=8'ha9;
	15'h21: q<=8'h00;
	15'h22: q<=8'h85;
	15'h23: q<=8'h01;
	15'h24: q<=8'h60;
	15'h25: q<=8'h20;
	15'h26: q<=8'h1b;
	15'h27: q<=8'h92;
	15'h28: q<=8'h20;
	15'h29: q<=8'hc5;
	15'h2a: q<=8'h92;
	15'h2b: q<=8'h20;
	15'h2c: q<=8'h8f;
	15'h2d: q<=8'h92;
	15'h2e: q<=8'h20;
	15'h2f: q<=8'h6f;
	15'h30: q<=8'h92;
	15'h31: q<=8'h20;
	15'h32: q<=8'h46;
	15'h33: q<=8'h92;
	15'h34: q<=8'h20;
	15'h35: q<=8'h9f;
	15'h36: q<=8'h92;
	15'h37: q<=8'h20;
	15'h38: q<=8'had;
	15'h39: q<=8'h92;
	15'h3a: q<=8'h20;
	15'h3b: q<=8'h6e;
	15'h3c: q<=8'hc1;
	15'h3d: q<=8'ha9;
	15'h3e: q<=8'hff;
	15'h3f: q<=8'h8d;
	15'h40: q<=8'h24;
	15'h41: q<=8'h01;
	15'h42: q<=8'h8d;
	15'h43: q<=8'h48;
	15'h44: q<=8'h01;
	15'h45: q<=8'ha9;
	15'h46: q<=8'h00;
	15'h47: q<=8'h8d;
	15'h48: q<=8'h23;
	15'h49: q<=8'h01;
	15'h4a: q<=8'h60;
	15'h4b: q<=8'ha9;
	15'h4c: q<=8'h10;
	15'h4d: q<=8'h8d;
	15'h4e: q<=8'h02;
	15'h4f: q<=8'h02;
	15'h50: q<=8'ha9;
	15'h51: q<=8'h00;
	15'h52: q<=8'h85;
	15'h53: q<=8'h29;
	15'h54: q<=8'h85;
	15'h55: q<=8'h2b;
	15'h56: q<=8'had;
	15'h57: q<=8'h21;
	15'h58: q<=8'h01;
	15'h59: q<=8'h85;
	15'h5a: q<=8'h2a;
	15'h5b: q<=8'h10;
	15'h5c: q<=8'h02;
	15'h5d: q<=8'hc6;
	15'h5e: q<=8'h2b;
	15'h5f: q<=8'ha2;
	15'h60: q<=8'h01;
	15'h61: q<=8'ha5;
	15'h62: q<=8'h2a;
	15'h63: q<=8'h0a;
	15'h64: q<=8'h66;
	15'h65: q<=8'h2a;
	15'h66: q<=8'h66;
	15'h67: q<=8'h29;
	15'h68: q<=8'hca;
	15'h69: q<=8'h10;
	15'h6a: q<=8'hf6;
	15'h6b: q<=8'ha5;
	15'h6c: q<=8'h29;
	15'h6d: q<=8'h18;
	15'h6e: q<=8'h6d;
	15'h6f: q<=8'h22;
	15'h70: q<=8'h01;
	15'h71: q<=8'h8d;
	15'h72: q<=8'h22;
	15'h73: q<=8'h01;
	15'h74: q<=8'ha5;
	15'h75: q<=8'h2a;
	15'h76: q<=8'h65;
	15'h77: q<=8'h68;
	15'h78: q<=8'h85;
	15'h79: q<=8'h68;
	15'h7a: q<=8'ha5;
	15'h7b: q<=8'h2b;
	15'h7c: q<=8'h65;
	15'h7d: q<=8'h69;
	15'h7e: q<=8'h85;
	15'h7f: q<=8'h69;
	15'h80: q<=8'ha5;
	15'h81: q<=8'h5f;
	15'h82: q<=8'h18;
	15'h83: q<=8'h69;
	15'h84: q<=8'h18;
	15'h85: q<=8'h85;
	15'h86: q<=8'h5f;
	15'h87: q<=8'ha5;
	15'h88: q<=8'h5b;
	15'h89: q<=8'h69;
	15'h8a: q<=8'h00;
	15'h8b: q<=8'h85;
	15'h8c: q<=8'h5b;
	15'h8d: q<=8'hc9;
	15'h8e: q<=8'hfc;
	15'h8f: q<=8'h90;
	15'h90: q<=8'h05;
	15'h91: q<=8'ha9;
	15'h92: q<=8'h01;
	15'h93: q<=8'h8d;
	15'h94: q<=8'h15;
	15'h95: q<=8'h01;
	15'h96: q<=8'ha5;
	15'h97: q<=8'h5f;
	15'h98: q<=8'h38;
	15'h99: q<=8'he5;
	15'h9a: q<=8'h5d;
	15'h9b: q<=8'ha5;
	15'h9c: q<=8'h5b;
	15'h9d: q<=8'hf0;
	15'h9e: q<=8'h02;
	15'h9f: q<=8'he9;
	15'ha0: q<=8'hff;
	15'ha1: q<=8'hd0;
	15'ha2: q<=8'h19;
	15'ha3: q<=8'ha5;
	15'ha4: q<=8'h5d;
	15'ha5: q<=8'h85;
	15'ha6: q<=8'h5f;
	15'ha7: q<=8'ha9;
	15'ha8: q<=8'hff;
	15'ha9: q<=8'h85;
	15'haa: q<=8'h5b;
	15'hab: q<=8'ha9;
	15'hac: q<=8'h04;
	15'had: q<=8'h24;
	15'hae: q<=8'h05;
	15'haf: q<=8'h30;
	15'hb0: q<=8'h02;
	15'hb1: q<=8'ha9;
	15'hb2: q<=8'h08;
	15'hb3: q<=8'h85;
	15'hb4: q<=8'h00;
	15'hb5: q<=8'ha6;
	15'hb6: q<=8'h3d;
	15'hb7: q<=8'ha9;
	15'hb8: q<=8'h00;
	15'hb9: q<=8'h9d;
	15'hba: q<=8'h02;
	15'hbb: q<=8'h01;
	15'hbc: q<=8'ha9;
	15'hbd: q<=8'hff;
	15'hbe: q<=8'h8d;
	15'hbf: q<=8'h14;
	15'hc0: q<=8'h01;
	15'hc1: q<=8'h4c;
	15'hc2: q<=8'h49;
	15'hc3: q<=8'h97;
	15'hc4: q<=8'had;
	15'hc5: q<=8'h26;
	15'hc6: q<=8'h01;
	15'hc7: q<=8'ha2;
	15'hc8: q<=8'h1c;
	15'hc9: q<=8'hca;
	15'hca: q<=8'hdd;
	15'hcb: q<=8'hfe;
	15'hcc: q<=8'h91;
	15'hcd: q<=8'h90;
	15'hce: q<=8'hfa;
	15'hcf: q<=8'ha0;
	15'hd0: q<=8'h04;
	15'hd1: q<=8'had;
	15'hd2: q<=8'h6a;
	15'hd3: q<=8'h01;
	15'hd4: q<=8'h29;
	15'hd5: q<=8'h04;
	15'hd6: q<=8'hf0;
	15'hd7: q<=8'h12;
	15'hd8: q<=8'had;
	15'hd9: q<=8'h1d;
	15'hda: q<=8'h07;
	15'hdb: q<=8'hc9;
	15'hdc: q<=8'h30;
	15'hdd: q<=8'h90;
	15'hde: q<=8'h01;
	15'hdf: q<=8'hc8;
	15'he0: q<=8'hc9;
	15'he1: q<=8'h50;
	15'he2: q<=8'h90;
	15'he3: q<=8'h01;
	15'he4: q<=8'hc8;
	15'he5: q<=8'hc9;
	15'he6: q<=8'h70;
	15'he7: q<=8'h90;
	15'he8: q<=8'h01;
	15'he9: q<=8'hc8;
	15'hea: q<=8'ha5;
	15'heb: q<=8'h09;
	15'hec: q<=8'h29;
	15'hed: q<=8'h43;
	15'hee: q<=8'hc9;
	15'hef: q<=8'h40;
	15'hf0: q<=8'hd0;
	15'hf1: q<=8'h02;
	15'hf2: q<=8'ha0;
	15'hf3: q<=8'h1b;
	15'hf4: q<=8'h84;
	15'hf5: q<=8'h29;
	15'hf6: q<=8'he4;
	15'hf7: q<=8'h29;
	15'hf8: q<=8'hb0;
	15'hf9: q<=8'h02;
	15'hfa: q<=8'ha6;
	15'hfb: q<=8'h29;
	15'hfc: q<=8'h8e;
	15'hfd: q<=8'h27;
	15'hfe: q<=8'h01;
	15'hff: q<=8'ha5;
	15'h100: q<=8'h05;
	15'h101: q<=8'h10;
	15'h102: q<=8'h05;
	15'h103: q<=8'ha9;
	15'h104: q<=8'h00;
	15'h105: q<=8'h8d;
	15'h106: q<=8'h26;
	15'h107: q<=8'h01;
	15'h108: q<=8'ha6;
	15'h109: q<=8'h3f;
	15'h10a: q<=8'h86;
	15'h10b: q<=8'h3d;
	15'h10c: q<=8'hf0;
	15'h10d: q<=8'h03;
	15'h10e: q<=8'h20;
	15'h10f: q<=8'hb2;
	15'h110: q<=8'h92;
	15'h111: q<=8'ha9;
	15'h112: q<=8'h04;
	15'h113: q<=8'h85;
	15'h114: q<=8'h7c;
	15'h115: q<=8'ha9;
	15'h116: q<=8'hff;
	15'h117: q<=8'h85;
	15'h118: q<=8'h5b;
	15'h119: q<=8'ha9;
	15'h11a: q<=8'h00;
	15'h11b: q<=8'h8d;
	15'h11c: q<=8'h00;
	15'h11d: q<=8'h02;
	15'h11e: q<=8'h85;
	15'h11f: q<=8'h51;
	15'h120: q<=8'h85;
	15'h121: q<=8'h7b;
	15'h122: q<=8'h8d;
	15'h123: q<=8'h05;
	15'h124: q<=8'h06;
	15'h125: q<=8'ha6;
	15'h126: q<=8'h05;
	15'h127: q<=8'h10;
	15'h128: q<=8'h1b;
	15'h129: q<=8'ha9;
	15'h12a: q<=8'h14;
	15'h12b: q<=8'h8d;
	15'h12c: q<=8'h05;
	15'h12d: q<=8'h06;
	15'h12e: q<=8'ha9;
	15'h12f: q<=8'hff;
	15'h130: q<=8'h8d;
	15'h131: q<=8'h11;
	15'h132: q<=8'h01;
	15'h133: q<=8'ha9;
	15'h134: q<=8'h16;
	15'h135: q<=8'h85;
	15'h136: q<=8'h00;
	15'h137: q<=8'ha9;
	15'h138: q<=8'h08;
	15'h139: q<=8'h85;
	15'h13a: q<=8'h01;
	15'h13b: q<=8'ha9;
	15'h13c: q<=8'h00;
	15'h13d: q<=8'h85;
	15'h13e: q<=8'h9f;
	15'h13f: q<=8'h20;
	15'h140: q<=8'h96;
	15'h141: q<=8'hc1;
	15'h142: q<=8'ha9;
	15'h143: q<=8'h10;
	15'h144: q<=8'h85;
	15'h145: q<=8'h04;
	15'h146: q<=8'h20;
	15'h147: q<=8'had;
	15'h148: q<=8'h92;
	15'h149: q<=8'hce;
	15'h14a: q<=8'h05;
	15'h14b: q<=8'h06;
	15'h14c: q<=8'h10;
	15'h14d: q<=8'h1b;
	15'h14e: q<=8'hf8;
	15'h14f: q<=8'ha5;
	15'h150: q<=8'h04;
	15'h151: q<=8'h38;
	15'h152: q<=8'he9;
	15'h153: q<=8'h01;
	15'h154: q<=8'h85;
	15'h155: q<=8'h04;
	15'h156: q<=8'hd8;
	15'h157: q<=8'h10;
	15'h158: q<=8'h04;
	15'h159: q<=8'ha9;
	15'h15a: q<=8'h10;
	15'h15b: q<=8'h85;
	15'h15c: q<=8'h4e;
	15'h15d: q<=8'hc9;
	15'h15e: q<=8'h03;
	15'h15f: q<=8'hd0;
	15'h160: q<=8'h03;
	15'h161: q<=8'h20;
	15'h162: q<=8'hfe;
	15'h163: q<=8'hcc;
	15'h164: q<=8'ha9;
	15'h165: q<=8'h14;
	15'h166: q<=8'h8d;
	15'h167: q<=8'h05;
	15'h168: q<=8'h06;
	15'h169: q<=8'h20;
	15'h16a: q<=8'hab;
	15'h16b: q<=8'hb0;
	15'h16c: q<=8'ha9;
	15'h16d: q<=8'h18;
	15'h16e: q<=8'ha4;
	15'h16f: q<=8'h04;
	15'h170: q<=8'hc0;
	15'h171: q<=8'h08;
	15'h172: q<=8'hb0;
	15'h173: q<=8'h02;
	15'h174: q<=8'ha9;
	15'h175: q<=8'h78;
	15'h176: q<=8'h25;
	15'h177: q<=8'h4e;
	15'h178: q<=8'hf0;
	15'h179: q<=8'h34;
	15'h17a: q<=8'ha9;
	15'h17b: q<=8'h00;
	15'h17c: q<=8'h85;
	15'h17d: q<=8'h4e;
	15'h17e: q<=8'had;
	15'h17f: q<=8'h00;
	15'h180: q<=8'h02;
	15'h181: q<=8'ha8;
	15'h182: q<=8'ha6;
	15'h183: q<=8'h3d;
	15'h184: q<=8'h9d;
	15'h185: q<=8'h02;
	15'h186: q<=8'h01;
	15'h187: q<=8'hb9;
	15'h188: q<=8'hfe;
	15'h189: q<=8'h91;
	15'h18a: q<=8'h24;
	15'h18b: q<=8'h05;
	15'h18c: q<=8'h30;
	15'h18d: q<=8'h09;
	15'h18e: q<=8'ha0;
	15'h18f: q<=8'h01;
	15'h190: q<=8'h84;
	15'h191: q<=8'h48;
	15'h192: q<=8'had;
	15'h193: q<=8'hca;
	15'h194: q<=8'h60;
	15'h195: q<=8'h29;
	15'h196: q<=8'h07;
	15'h197: q<=8'h95;
	15'h198: q<=8'h46;
	15'h199: q<=8'h85;
	15'h19a: q<=8'h9f;
	15'h19b: q<=8'h20;
	15'h19c: q<=8'h96;
	15'h19d: q<=8'hc1;
	15'h19e: q<=8'h20;
	15'h19f: q<=8'hc5;
	15'h1a0: q<=8'h92;
	15'h1a1: q<=8'h20;
	15'h1a2: q<=8'h34;
	15'h1a3: q<=8'h92;
	15'h1a4: q<=8'h20;
	15'h1a5: q<=8'h31;
	15'h1a6: q<=8'ha8;
	15'h1a7: q<=8'ha9;
	15'h1a8: q<=8'h02;
	15'h1a9: q<=8'h85;
	15'h1aa: q<=8'h00;
	15'h1ab: q<=8'h20;
	15'h1ac: q<=8'had;
	15'h1ad: q<=8'h92;
	15'h1ae: q<=8'ha5;
	15'h1af: q<=8'h4e;
	15'h1b0: q<=8'h29;
	15'h1b1: q<=8'h07;
	15'h1b2: q<=8'h85;
	15'h1b3: q<=8'h4e;
	15'h1b4: q<=8'h60;
	15'h1b5: q<=8'h0a;
	15'h1b6: q<=8'haa;
	15'h1b7: q<=8'ha9;
	15'h1b8: q<=8'h00;
	15'h1b9: q<=8'h85;
	15'h1ba: q<=8'h29;
	15'h1bb: q<=8'hbd;
	15'h1bc: q<=8'hc6;
	15'h1bd: q<=8'h91;
	15'h1be: q<=8'h85;
	15'h1bf: q<=8'h2a;
	15'h1c0: q<=8'hbd;
	15'h1c1: q<=8'hc7;
	15'h1c2: q<=8'h91;
	15'h1c3: q<=8'h85;
	15'h1c4: q<=8'h2b;
	15'h1c5: q<=8'h60;
	15'h1c6: q<=8'h00;
	15'h1c7: q<=8'h00;
	15'h1c8: q<=8'h60;
	15'h1c9: q<=8'h00;
	15'h1ca: q<=8'h60;
	15'h1cb: q<=8'h01;
	15'h1cc: q<=8'h20;
	15'h1cd: q<=8'h03;
	15'h1ce: q<=8'h40;
	15'h1cf: q<=8'h05;
	15'h1d0: q<=8'h40;
	15'h1d1: q<=8'h07;
	15'h1d2: q<=8'h40;
	15'h1d3: q<=8'h09;
	15'h1d4: q<=8'h40;
	15'h1d5: q<=8'h11;
	15'h1d6: q<=8'h40;
	15'h1d7: q<=8'h13;
	15'h1d8: q<=8'h20;
	15'h1d9: q<=8'h15;
	15'h1da: q<=8'h00;
	15'h1db: q<=8'h17;
	15'h1dc: q<=8'h80;
	15'h1dd: q<=8'h18;
	15'h1de: q<=8'h80;
	15'h1df: q<=8'h20;
	15'h1e0: q<=8'h60;
	15'h1e1: q<=8'h22;
	15'h1e2: q<=8'h80;
	15'h1e3: q<=8'h24;
	15'h1e4: q<=8'h60;
	15'h1e5: q<=8'h26;
	15'h1e6: q<=8'h00;
	15'h1e7: q<=8'h30;
	15'h1e8: q<=8'h00;
	15'h1e9: q<=8'h34;
	15'h1ea: q<=8'h20;
	15'h1eb: q<=8'h38;
	15'h1ec: q<=8'h50;
	15'h1ed: q<=8'h41;
	15'h1ee: q<=8'h90;
	15'h1ef: q<=8'h43;
	15'h1f0: q<=8'h20;
	15'h1f1: q<=8'h47;
	15'h1f2: q<=8'h10;
	15'h1f3: q<=8'h53;
	15'h1f4: q<=8'h10;
	15'h1f5: q<=8'h58;
	15'h1f6: q<=8'h40;
	15'h1f7: q<=8'h62;
	15'h1f8: q<=8'h60;
	15'h1f9: q<=8'h65;
	15'h1fa: q<=8'h60;
	15'h1fb: q<=8'h76;
	15'h1fc: q<=8'h80;
	15'h1fd: q<=8'h89;
	15'h1fe: q<=8'h00;
	15'h1ff: q<=8'h02;
	15'h200: q<=8'h04;
	15'h201: q<=8'h06;
	15'h202: q<=8'h08;
	15'h203: q<=8'h0a;
	15'h204: q<=8'h0c;
	15'h205: q<=8'h0e;
	15'h206: q<=8'h10;
	15'h207: q<=8'h13;
	15'h208: q<=8'h15;
	15'h209: q<=8'h17;
	15'h20a: q<=8'h19;
	15'h20b: q<=8'h1b;
	15'h20c: q<=8'h1e;
	15'h20d: q<=8'h20;
	15'h20e: q<=8'h23;
	15'h20f: q<=8'h27;
	15'h210: q<=8'h2b;
	15'h211: q<=8'h2e;
	15'h212: q<=8'h30;
	15'h213: q<=8'h33;
	15'h214: q<=8'h37;
	15'h215: q<=8'h3b;
	15'h216: q<=8'h3e;
	15'h217: q<=8'h40;
	15'h218: q<=8'h48;
	15'h219: q<=8'h50;
	15'h21a: q<=8'hff;
	15'h21b: q<=8'ha9;
	15'h21c: q<=8'h0e;
	15'h21d: q<=8'h8d;
	15'h21e: q<=8'h00;
	15'h21f: q<=8'h02;
	15'h220: q<=8'ha9;
	15'h221: q<=8'hf0;
	15'h222: q<=8'h85;
	15'h223: q<=8'h51;
	15'h224: q<=8'ha9;
	15'h225: q<=8'h00;
	15'h226: q<=8'h8d;
	15'h227: q<=8'h06;
	15'h228: q<=8'h01;
	15'h229: q<=8'ha9;
	15'h22a: q<=8'h0f;
	15'h22b: q<=8'h8d;
	15'h22c: q<=8'h01;
	15'h22d: q<=8'h02;
	15'h22e: q<=8'ha9;
	15'h22f: q<=8'h10;
	15'h230: q<=8'h8d;
	15'h231: q<=8'h02;
	15'h232: q<=8'h02;
	15'h233: q<=8'h60;
	15'h234: q<=8'had;
	15'h235: q<=8'h5b;
	15'h236: q<=8'h01;
	15'h237: q<=8'h8d;
	15'h238: q<=8'hab;
	15'h239: q<=8'h03;
	15'h23a: q<=8'had;
	15'h23b: q<=8'h5a;
	15'h23c: q<=8'h01;
	15'h23d: q<=8'ha2;
	15'h23e: q<=8'h0f;
	15'h23f: q<=8'h9d;
	15'h240: q<=8'hac;
	15'h241: q<=8'h03;
	15'h242: q<=8'hca;
	15'h243: q<=8'h10;
	15'h244: q<=8'hfa;
	15'h245: q<=8'h60;
	15'h246: q<=8'ha9;
	15'h247: q<=8'h00;
	15'h248: q<=8'ha2;
	15'h249: q<=8'h3f;
	15'h24a: q<=8'h9d;
	15'h24b: q<=8'h43;
	15'h24c: q<=8'h02;
	15'h24d: q<=8'hca;
	15'h24e: q<=8'h10;
	15'h24f: q<=8'hfa;
	15'h250: q<=8'hae;
	15'h251: q<=8'hab;
	15'h252: q<=8'h03;
	15'h253: q<=8'hca;
	15'h254: q<=8'had;
	15'h255: q<=8'hca;
	15'h256: q<=8'h60;
	15'h257: q<=8'h29;
	15'h258: q<=8'h0f;
	15'h259: q<=8'h9d;
	15'h25a: q<=8'h03;
	15'h25b: q<=8'h02;
	15'h25c: q<=8'h8a;
	15'h25d: q<=8'h0a;
	15'h25e: q<=8'h0a;
	15'h25f: q<=8'h0a;
	15'h260: q<=8'h0a;
	15'h261: q<=8'h1d;
	15'h262: q<=8'h03;
	15'h263: q<=8'h02;
	15'h264: q<=8'hd0;
	15'h265: q<=8'h02;
	15'h266: q<=8'ha9;
	15'h267: q<=8'h0f;
	15'h268: q<=8'h9d;
	15'h269: q<=8'h43;
	15'h26a: q<=8'h02;
	15'h26b: q<=8'hca;
	15'h26c: q<=8'h10;
	15'h26d: q<=8'he6;
	15'h26e: q<=8'h60;
	15'h26f: q<=8'ha2;
	15'h270: q<=8'h06;
	15'h271: q<=8'ha9;
	15'h272: q<=8'h00;
	15'h273: q<=8'h9d;
	15'h274: q<=8'hdf;
	15'h275: q<=8'h02;
	15'h276: q<=8'hca;
	15'h277: q<=8'h10;
	15'h278: q<=8'hfa;
	15'h279: q<=8'h8d;
	15'h27a: q<=8'h08;
	15'h27b: q<=8'h01;
	15'h27c: q<=8'h8d;
	15'h27d: q<=8'h09;
	15'h27e: q<=8'h01;
	15'h27f: q<=8'h8d;
	15'h280: q<=8'h45;
	15'h281: q<=8'h01;
	15'h282: q<=8'h8d;
	15'h283: q<=8'h42;
	15'h284: q<=8'h01;
	15'h285: q<=8'h8d;
	15'h286: q<=8'h44;
	15'h287: q<=8'h01;
	15'h288: q<=8'h8d;
	15'h289: q<=8'h43;
	15'h28a: q<=8'h01;
	15'h28b: q<=8'h8d;
	15'h28c: q<=8'h46;
	15'h28d: q<=8'h01;
	15'h28e: q<=8'h60;
	15'h28f: q<=8'ha9;
	15'h290: q<=8'h00;
	15'h291: q<=8'ha2;
	15'h292: q<=8'h0b;
	15'h293: q<=8'h9d;
	15'h294: q<=8'hd3;
	15'h295: q<=8'h02;
	15'h296: q<=8'hca;
	15'h297: q<=8'h10;
	15'h298: q<=8'hfa;
	15'h299: q<=8'h8d;
	15'h29a: q<=8'h35;
	15'h29b: q<=8'h01;
	15'h29c: q<=8'h85;
	15'h29d: q<=8'ha6;
	15'h29e: q<=8'h60;
	15'h29f: q<=8'ha2;
	15'h2a0: q<=8'h07;
	15'h2a1: q<=8'ha9;
	15'h2a2: q<=8'h00;
	15'h2a3: q<=8'h9d;
	15'h2a4: q<=8'h0a;
	15'h2a5: q<=8'h03;
	15'h2a6: q<=8'hca;
	15'h2a7: q<=8'h10;
	15'h2a8: q<=8'hfa;
	15'h2a9: q<=8'h8d;
	15'h2aa: q<=8'h16;
	15'h2ab: q<=8'h01;
	15'h2ac: q<=8'h60;
	15'h2ad: q<=8'ha9;
	15'h2ae: q<=8'h00;
	15'h2af: q<=8'h85;
	15'h2b0: q<=8'h50;
	15'h2b1: q<=8'h60;
	15'h2b2: q<=8'ha2;
	15'h2b3: q<=8'h11;
	15'h2b4: q<=8'hbd;
	15'h2b5: q<=8'haa;
	15'h2b6: q<=8'h03;
	15'h2b7: q<=8'hbc;
	15'h2b8: q<=8'hbc;
	15'h2b9: q<=8'h03;
	15'h2ba: q<=8'h9d;
	15'h2bb: q<=8'hbc;
	15'h2bc: q<=8'h03;
	15'h2bd: q<=8'h98;
	15'h2be: q<=8'h9d;
	15'h2bf: q<=8'haa;
	15'h2c0: q<=8'h03;
	15'h2c1: q<=8'hca;
	15'h2c2: q<=8'h10;
	15'h2c3: q<=8'hf0;
	15'h2c4: q<=8'h60;
	15'h2c5: q<=8'ha5;
	15'h2c6: q<=8'h9f;
	15'h2c7: q<=8'hc9;
	15'h2c8: q<=8'h62;
	15'h2c9: q<=8'h90;
	15'h2ca: q<=8'h07;
	15'h2cb: q<=8'had;
	15'h2cc: q<=8'hda;
	15'h2cd: q<=8'h60;
	15'h2ce: q<=8'h29;
	15'h2cf: q<=8'h1f;
	15'h2d0: q<=8'h09;
	15'h2d1: q<=8'h40;
	15'h2d2: q<=8'h85;
	15'h2d3: q<=8'h2b;
	15'h2d4: q<=8'he6;
	15'h2d5: q<=8'h2b;
	15'h2d6: q<=8'ha2;
	15'h2d7: q<=8'h6f;
	15'h2d8: q<=8'h86;
	15'h2d9: q<=8'h37;
	15'h2da: q<=8'ha6;
	15'h2db: q<=8'h37;
	15'h2dc: q<=8'hbd;
	15'h2dd: q<=8'h07;
	15'h2de: q<=8'h96;
	15'h2df: q<=8'h85;
	15'h2e0: q<=8'h3c;
	15'h2e1: q<=8'hbd;
	15'h2e2: q<=8'h06;
	15'h2e3: q<=8'h96;
	15'h2e4: q<=8'h85;
	15'h2e5: q<=8'h3b;
	15'h2e6: q<=8'hbd;
	15'h2e7: q<=8'h05;
	15'h2e8: q<=8'h96;
	15'h2e9: q<=8'h85;
	15'h2ea: q<=8'h2d;
	15'h2eb: q<=8'hbd;
	15'h2ec: q<=8'h04;
	15'h2ed: q<=8'h96;
	15'h2ee: q<=8'h85;
	15'h2ef: q<=8'h2c;
	15'h2f0: q<=8'ha9;
	15'h2f1: q<=8'h01;
	15'h2f2: q<=8'h85;
	15'h2f3: q<=8'h38;
	15'h2f4: q<=8'ha0;
	15'h2f5: q<=8'h00;
	15'h2f6: q<=8'hb1;
	15'h2f7: q<=8'h2c;
	15'h2f8: q<=8'h8d;
	15'h2f9: q<=8'h5e;
	15'h2fa: q<=8'h01;
	15'h2fb: q<=8'hf0;
	15'h2fc: q<=8'h1c;
	15'h2fd: q<=8'ha5;
	15'h2fe: q<=8'h2b;
	15'h2ff: q<=8'hc8;
	15'h300: q<=8'hd1;
	15'h301: q<=8'h2c;
	15'h302: q<=8'hc8;
	15'h303: q<=8'h90;
	15'h304: q<=8'h0e;
	15'h305: q<=8'hd1;
	15'h306: q<=8'h2c;
	15'h307: q<=8'hd0;
	15'h308: q<=8'h01;
	15'h309: q<=8'h18;
	15'h30a: q<=8'hb0;
	15'h30b: q<=8'h07;
	15'h30c: q<=8'hc8;
	15'h30d: q<=8'h20;
	15'h30e: q<=8'h77;
	15'h30f: q<=8'h96;
	15'h310: q<=8'h4c;
	15'h311: q<=8'h19;
	15'h312: q<=8'h93;
	15'h313: q<=8'h20;
	15'h314: q<=8'h83;
	15'h315: q<=8'h96;
	15'h316: q<=8'h18;
	15'h317: q<=8'h90;
	15'h318: q<=8'hdd;
	15'h319: q<=8'ha0;
	15'h31a: q<=8'h00;
	15'h31b: q<=8'h91;
	15'h31c: q<=8'h3b;
	15'h31d: q<=8'ha5;
	15'h31e: q<=8'h37;
	15'h31f: q<=8'h38;
	15'h320: q<=8'he9;
	15'h321: q<=8'h04;
	15'h322: q<=8'h85;
	15'h323: q<=8'h37;
	15'h324: q<=8'hc9;
	15'h325: q<=8'hff;
	15'h326: q<=8'hd0;
	15'h327: q<=8'hb2;
	15'h328: q<=8'had;
	15'h329: q<=8'h6a;
	15'h32a: q<=8'h01;
	15'h32b: q<=8'h29;
	15'h32c: q<=8'h03;
	15'h32d: q<=8'hc9;
	15'h32e: q<=8'h01;
	15'h32f: q<=8'hd0;
	15'h330: q<=8'h1c;
	15'h331: q<=8'hce;
	15'h332: q<=8'h1a;
	15'h333: q<=8'h01;
	15'h334: q<=8'had;
	15'h335: q<=8'h60;
	15'h336: q<=8'h01;
	15'h337: q<=8'h49;
	15'h338: q<=8'hff;
	15'h339: q<=8'h4a;
	15'h33a: q<=8'h4a;
	15'h33b: q<=8'h4a;
	15'h33c: q<=8'h6d;
	15'h33d: q<=8'h60;
	15'h33e: q<=8'h01;
	15'h33f: q<=8'h8d;
	15'h340: q<=8'h60;
	15'h341: q<=8'h01;
	15'h342: q<=8'ha5;
	15'h343: q<=8'h9f;
	15'h344: q<=8'hc9;
	15'h345: q<=8'h11;
	15'h346: q<=8'hb0;
	15'h347: q<=8'h02;
	15'h348: q<=8'hc6;
	15'h349: q<=8'hb3;
	15'h34a: q<=8'hb8;
	15'h34b: q<=8'h50;
	15'h34c: q<=8'h35;
	15'h34d: q<=8'hc9;
	15'h34e: q<=8'h02;
	15'h34f: q<=8'hd0;
	15'h350: q<=8'h31;
	15'h351: q<=8'hee;
	15'h352: q<=8'h1a;
	15'h353: q<=8'h01;
	15'h354: q<=8'had;
	15'h355: q<=8'h1a;
	15'h356: q<=8'h01;
	15'h357: q<=8'hc9;
	15'h358: q<=8'h03;
	15'h359: q<=8'h90;
	15'h35a: q<=8'h05;
	15'h35b: q<=8'ha9;
	15'h35c: q<=8'h03;
	15'h35d: q<=8'h8d;
	15'h35e: q<=8'h1a;
	15'h35f: q<=8'h01;
	15'h360: q<=8'had;
	15'h361: q<=8'h60;
	15'h362: q<=8'h01;
	15'h363: q<=8'h4a;
	15'h364: q<=8'h4a;
	15'h365: q<=8'h4a;
	15'h366: q<=8'h09;
	15'h367: q<=8'he0;
	15'h368: q<=8'h6d;
	15'h369: q<=8'h60;
	15'h36a: q<=8'h01;
	15'h36b: q<=8'h8d;
	15'h36c: q<=8'h60;
	15'h36d: q<=8'h01;
	15'h36e: q<=8'had;
	15'h36f: q<=8'h5b;
	15'h370: q<=8'h01;
	15'h371: q<=8'h4a;
	15'h372: q<=8'h4a;
	15'h373: q<=8'h4a;
	15'h374: q<=8'h6d;
	15'h375: q<=8'h5b;
	15'h376: q<=8'h01;
	15'h377: q<=8'h8d;
	15'h378: q<=8'h5b;
	15'h379: q<=8'h01;
	15'h37a: q<=8'had;
	15'h37b: q<=8'h6d;
	15'h37c: q<=8'h01;
	15'h37d: q<=8'h09;
	15'h37e: q<=8'h40;
	15'h37f: q<=8'h8d;
	15'h380: q<=8'h6d;
	15'h381: q<=8'h01;
	15'h382: q<=8'had;
	15'h383: q<=8'h63;
	15'h384: q<=8'h01;
	15'h385: q<=8'h20;
	15'h386: q<=8'he0;
	15'h387: q<=8'h93;
	15'h388: q<=8'h8d;
	15'h389: q<=8'h63;
	15'h38a: q<=8'h01;
	15'h38b: q<=8'h8c;
	15'h38c: q<=8'h68;
	15'h38d: q<=8'h01;
	15'h38e: q<=8'h8e;
	15'h38f: q<=8'h54;
	15'h390: q<=8'h01;
	15'h391: q<=8'had;
	15'h392: q<=8'h20;
	15'h393: q<=8'h01;
	15'h394: q<=8'h20;
	15'h395: q<=8'he0;
	15'h396: q<=8'h93;
	15'h397: q<=8'h8d;
	15'h398: q<=8'h20;
	15'h399: q<=8'h01;
	15'h39a: q<=8'h8c;
	15'h39b: q<=8'h18;
	15'h39c: q<=8'h01;
	15'h39d: q<=8'h86;
	15'h39e: q<=8'ha7;
	15'h39f: q<=8'had;
	15'h3a0: q<=8'h60;
	15'h3a1: q<=8'h01;
	15'h3a2: q<=8'h20;
	15'h3a3: q<=8'he0;
	15'h3a4: q<=8'h93;
	15'h3a5: q<=8'h8d;
	15'h3a6: q<=8'h60;
	15'h3a7: q<=8'h01;
	15'h3a8: q<=8'h8d;
	15'h3a9: q<=8'h62;
	15'h3aa: q<=8'h01;
	15'h3ab: q<=8'h8c;
	15'h3ac: q<=8'h67;
	15'h3ad: q<=8'h01;
	15'h3ae: q<=8'h8c;
	15'h3af: q<=8'h65;
	15'h3b0: q<=8'h01;
	15'h3b1: q<=8'h8e;
	15'h3b2: q<=8'h51;
	15'h3b3: q<=8'h01;
	15'h3b4: q<=8'h8e;
	15'h3b5: q<=8'h53;
	15'h3b6: q<=8'h01;
	15'h3b7: q<=8'h8e;
	15'h3b8: q<=8'h52;
	15'h3b9: q<=8'h01;
	15'h3ba: q<=8'had;
	15'h3bb: q<=8'h60;
	15'h3bc: q<=8'h01;
	15'h3bd: q<=8'h0a;
	15'h3be: q<=8'h8d;
	15'h3bf: q<=8'h64;
	15'h3c0: q<=8'h01;
	15'h3c1: q<=8'had;
	15'h3c2: q<=8'h65;
	15'h3c3: q<=8'h01;
	15'h3c4: q<=8'h2a;
	15'h3c5: q<=8'h8d;
	15'h3c6: q<=8'h69;
	15'h3c7: q<=8'h01;
	15'h3c8: q<=8'ha9;
	15'h3c9: q<=8'h06;
	15'h3ca: q<=8'h8d;
	15'h3cb: q<=8'h55;
	15'h3cc: q<=8'h01;
	15'h3cd: q<=8'ha9;
	15'h3ce: q<=8'ha0;
	15'h3cf: q<=8'h8d;
	15'h3d0: q<=8'h61;
	15'h3d1: q<=8'h01;
	15'h3d2: q<=8'ha9;
	15'h3d3: q<=8'hfe;
	15'h3d4: q<=8'h8d;
	15'h3d5: q<=8'h66;
	15'h3d6: q<=8'h01;
	15'h3d7: q<=8'ha9;
	15'h3d8: q<=8'h01;
	15'h3d9: q<=8'h8d;
	15'h3da: q<=8'h4a;
	15'h3db: q<=8'h01;
	15'h3dc: q<=8'h8d;
	15'h3dd: q<=8'h49;
	15'h3de: q<=8'h01;
	15'h3df: q<=8'h60;
	15'h3e0: q<=8'ha0;
	15'h3e1: q<=8'hff;
	15'h3e2: q<=8'h84;
	15'h3e3: q<=8'h29;
	15'h3e4: q<=8'h0a;
	15'h3e5: q<=8'h26;
	15'h3e6: q<=8'h29;
	15'h3e7: q<=8'h0a;
	15'h3e8: q<=8'h26;
	15'h3e9: q<=8'h29;
	15'h3ea: q<=8'h0a;
	15'h3eb: q<=8'h26;
	15'h3ec: q<=8'h29;
	15'h3ed: q<=8'ha4;
	15'h3ee: q<=8'h29;
	15'h3ef: q<=8'h48;
	15'h3f0: q<=8'h98;
	15'h3f1: q<=8'h49;
	15'h3f2: q<=8'hff;
	15'h3f3: q<=8'h18;
	15'h3f4: q<=8'h69;
	15'h3f5: q<=8'h0d;
	15'h3f6: q<=8'h4a;
	15'h3f7: q<=8'haa;
	15'h3f8: q<=8'h68;
	15'h3f9: q<=8'h60;
	15'h3fa: q<=8'h08;
	15'h3fb: q<=8'h01;
	15'h3fc: q<=8'h14;
	15'h3fd: q<=8'h50;
	15'h3fe: q<=8'hfd;
	15'h3ff: q<=8'h02;
	15'h400: q<=8'h15;
	15'h401: q<=8'h40;
	15'h402: q<=8'h14;
	15'h403: q<=8'h02;
	15'h404: q<=8'h41;
	15'h405: q<=8'h63;
	15'h406: q<=8'h0a;
	15'h407: q<=8'h04;
	15'h408: q<=8'h01;
	15'h409: q<=8'h09;
	15'h40a: q<=8'h01;
	15'h40b: q<=8'h01;
	15'h40c: q<=8'h01;
	15'h40d: q<=8'h02;
	15'h40e: q<=8'h03;
	15'h40f: q<=8'h02;
	15'h410: q<=8'h02;
	15'h411: q<=8'h03;
	15'h412: q<=8'h03;
	15'h413: q<=8'h02;
	15'h414: q<=8'h0a;
	15'h415: q<=8'h40;
	15'h416: q<=8'h02;
	15'h417: q<=8'h02;
	15'h418: q<=8'h41;
	15'h419: q<=8'h63;
	15'h41a: q<=8'h03;
	15'h41b: q<=8'h08;
	15'h41c: q<=8'h01;
	15'h41d: q<=8'h08;
	15'h41e: q<=8'hd4;
	15'h41f: q<=8'hfb;
	15'h420: q<=8'h04;
	15'h421: q<=8'h09;
	15'h422: q<=8'h10;
	15'h423: q<=8'haf;
	15'h424: q<=8'hac;
	15'h425: q<=8'hac;
	15'h426: q<=8'hac;
	15'h427: q<=8'ha8;
	15'h428: q<=8'ha4;
	15'h429: q<=8'ha0;
	15'h42a: q<=8'ha0;
	15'h42b: q<=8'h08;
	15'h42c: q<=8'h11;
	15'h42d: q<=8'h19;
	15'h42e: q<=8'haf;
	15'h42f: q<=8'hfd;
	15'h430: q<=8'h08;
	15'h431: q<=8'h1a;
	15'h432: q<=8'h20;
	15'h433: q<=8'h9d;
	15'h434: q<=8'hfd;
	15'h435: q<=8'h08;
	15'h436: q<=8'h21;
	15'h437: q<=8'h27;
	15'h438: q<=8'h94;
	15'h439: q<=8'hfd;
	15'h43a: q<=8'h08;
	15'h43b: q<=8'h28;
	15'h43c: q<=8'h30;
	15'h43d: q<=8'h92;
	15'h43e: q<=8'hff;
	15'h43f: q<=8'h08;
	15'h440: q<=8'h31;
	15'h441: q<=8'h40;
	15'h442: q<=8'h88;
	15'h443: q<=8'hff;
	15'h444: q<=8'h0c;
	15'h445: q<=8'h41;
	15'h446: q<=8'h63;
	15'h447: q<=8'h60;
	15'h448: q<=8'h41;
	15'h449: q<=8'h0a;
	15'h44a: q<=8'h01;
	15'h44b: q<=8'h63;
	15'h44c: q<=8'hc0;
	15'h44d: q<=8'h0a;
	15'h44e: q<=8'h01;
	15'h44f: q<=8'h14;
	15'h450: q<=8'h00;
	15'h451: q<=8'h0a;
	15'h452: q<=8'h15;
	15'h453: q<=8'h20;
	15'h454: q<=8'hd0;
	15'h455: q<=8'h0a;
	15'h456: q<=8'h21;
	15'h457: q<=8'h30;
	15'h458: q<=8'hd8;
	15'h459: q<=8'h0a;
	15'h45a: q<=8'h31;
	15'h45b: q<=8'h63;
	15'h45c: q<=8'hd0;
	15'h45d: q<=8'h02;
	15'h45e: q<=8'h01;
	15'h45f: q<=8'h20;
	15'h460: q<=8'ha0;
	15'h461: q<=8'h02;
	15'h462: q<=8'h21;
	15'h463: q<=8'h40;
	15'h464: q<=8'ha0;
	15'h465: q<=8'h02;
	15'h466: q<=8'h41;
	15'h467: q<=8'h63;
	15'h468: q<=8'hc0;
	15'h469: q<=8'h02;
	15'h46a: q<=8'h01;
	15'h46b: q<=8'h30;
	15'h46c: q<=8'h04;
	15'h46d: q<=8'h02;
	15'h46e: q<=8'h31;
	15'h46f: q<=8'h40;
	15'h470: q<=8'h06;
	15'h471: q<=8'h02;
	15'h472: q<=8'h41;
	15'h473: q<=8'h63;
	15'h474: q<=8'h08;
	15'h475: q<=8'h02;
	15'h476: q<=8'h01;
	15'h477: q<=8'h20;
	15'h478: q<=8'h01;
	15'h479: q<=8'h02;
	15'h47a: q<=8'h21;
	15'h47b: q<=8'h28;
	15'h47c: q<=8'h03;
	15'h47d: q<=8'h02;
	15'h47e: q<=8'h29;
	15'h47f: q<=8'h63;
	15'h480: q<=8'h02;
	15'h481: q<=8'h02;
	15'h482: q<=8'h01;
	15'h483: q<=8'h30;
	15'h484: q<=8'h01;
	15'h485: q<=8'h02;
	15'h486: q<=8'h31;
	15'h487: q<=8'h63;
	15'h488: q<=8'h03;
	15'h489: q<=8'h04;
	15'h48a: q<=8'h01;
	15'h48b: q<=8'h04;
	15'h48c: q<=8'h00;
	15'h48d: q<=8'h00;
	15'h48e: q<=8'h00;
	15'h48f: q<=8'h01;
	15'h490: q<=8'h02;
	15'h491: q<=8'h05;
	15'h492: q<=8'h10;
	15'h493: q<=8'h02;
	15'h494: q<=8'h02;
	15'h495: q<=8'h11;
	15'h496: q<=8'h13;
	15'h497: q<=8'h00;
	15'h498: q<=8'h02;
	15'h499: q<=8'h14;
	15'h49a: q<=8'h20;
	15'h49b: q<=8'h01;
	15'h49c: q<=8'h02;
	15'h49d: q<=8'h23;
	15'h49e: q<=8'h27;
	15'h49f: q<=8'h01;
	15'h4a0: q<=8'h02;
	15'h4a1: q<=8'h2c;
	15'h4a2: q<=8'h63;
	15'h4a3: q<=8'h01;
	15'h4a4: q<=8'h00;
	15'h4a5: q<=8'h04;
	15'h4a6: q<=8'h01;
	15'h4a7: q<=8'h06;
	15'h4a8: q<=8'h00;
	15'h4a9: q<=8'h00;
	15'h4aa: q<=8'h00;
	15'h4ab: q<=8'h02;
	15'h4ac: q<=8'h03;
	15'h4ad: q<=8'h04;
	15'h4ae: q<=8'h02;
	15'h4af: q<=8'h07;
	15'h4b0: q<=8'h0a;
	15'h4b1: q<=8'h04;
	15'h4b2: q<=8'h02;
	15'h4b3: q<=8'h0b;
	15'h4b4: q<=8'h10;
	15'h4b5: q<=8'h03;
	15'h4b6: q<=8'h02;
	15'h4b7: q<=8'h14;
	15'h4b8: q<=8'h19;
	15'h4b9: q<=8'h02;
	15'h4ba: q<=8'h04;
	15'h4bb: q<=8'h1a;
	15'h4bc: q<=8'h20;
	15'h4bd: q<=8'h01;
	15'h4be: q<=8'h02;
	15'h4bf: q<=8'h02;
	15'h4c0: q<=8'h02;
	15'h4c1: q<=8'h01;
	15'h4c2: q<=8'h01;
	15'h4c3: q<=8'h02;
	15'h4c4: q<=8'h02;
	15'h4c5: q<=8'h35;
	15'h4c6: q<=8'h27;
	15'h4c7: q<=8'h01;
	15'h4c8: q<=8'h02;
	15'h4c9: q<=8'h2b;
	15'h4ca: q<=8'h63;
	15'h4cb: q<=8'h01;
	15'h4cc: q<=8'h00;
	15'h4cd: q<=8'h02;
	15'h4ce: q<=8'h01;
	15'h4cf: q<=8'h04;
	15'h4d0: q<=8'h01;
	15'h4d1: q<=8'h02;
	15'h4d2: q<=8'h05;
	15'h4d3: q<=8'h63;
	15'h4d4: q<=8'h00;
	15'h4d5: q<=8'h00;
	15'h4d6: q<=8'h02;
	15'h4d7: q<=8'h01;
	15'h4d8: q<=8'h04;
	15'h4d9: q<=8'h04;
	15'h4da: q<=8'h02;
	15'h4db: q<=8'h05;
	15'h4dc: q<=8'h10;
	15'h4dd: q<=8'h05;
	15'h4de: q<=8'h02;
	15'h4df: q<=8'h11;
	15'h4e0: q<=8'h13;
	15'h4e1: q<=8'h03;
	15'h4e2: q<=8'h02;
	15'h4e3: q<=8'h14;
	15'h4e4: q<=8'h19;
	15'h4e5: q<=8'h04;
	15'h4e6: q<=8'h02;
	15'h4e7: q<=8'h1a;
	15'h4e8: q<=8'h63;
	15'h4e9: q<=8'h05;
	15'h4ea: q<=8'h00;
	15'h4eb: q<=8'h04;
	15'h4ec: q<=8'h01;
	15'h4ed: q<=8'h04;
	15'h4ee: q<=8'h00;
	15'h4ef: q<=8'h00;
	15'h4f0: q<=8'h01;
	15'h4f1: q<=8'h00;
	15'h4f2: q<=8'h02;
	15'h4f3: q<=8'h05;
	15'h4f4: q<=8'h10;
	15'h4f5: q<=8'h01;
	15'h4f6: q<=8'h02;
	15'h4f7: q<=8'h11;
	15'h4f8: q<=8'h20;
	15'h4f9: q<=8'h01;
	15'h4fa: q<=8'h02;
	15'h4fb: q<=8'h21;
	15'h4fc: q<=8'h27;
	15'h4fd: q<=8'h01;
	15'h4fe: q<=8'h02;
	15'h4ff: q<=8'h28;
	15'h500: q<=8'h63;
	15'h501: q<=8'h01;
	15'h502: q<=8'h00;
	15'h503: q<=8'h04;
	15'h504: q<=8'h01;
	15'h505: q<=8'h05;
	15'h506: q<=8'h00;
	15'h507: q<=8'h00;
	15'h508: q<=8'h01;
	15'h509: q<=8'h00;
	15'h50a: q<=8'h01;
	15'h50b: q<=8'h02;
	15'h50c: q<=8'h06;
	15'h50d: q<=8'h10;
	15'h50e: q<=8'h02;
	15'h50f: q<=8'h02;
	15'h510: q<=8'h11;
	15'h511: q<=8'h1a;
	15'h512: q<=8'h01;
	15'h513: q<=8'h02;
	15'h514: q<=8'h1b;
	15'h515: q<=8'h20;
	15'h516: q<=8'h01;
	15'h517: q<=8'h02;
	15'h518: q<=8'h21;
	15'h519: q<=8'h2c;
	15'h51a: q<=8'h02;
	15'h51b: q<=8'h02;
	15'h51c: q<=8'h2d;
	15'h51d: q<=8'h63;
	15'h51e: q<=8'h03;
	15'h51f: q<=8'h00;
	15'h520: q<=8'h02;
	15'h521: q<=8'h11;
	15'h522: q<=8'h20;
	15'h523: q<=8'h02;
	15'h524: q<=8'h02;
	15'h525: q<=8'h21;
	15'h526: q<=8'h63;
	15'h527: q<=8'h01;
	15'h528: q<=8'h00;
	15'h529: q<=8'h04;
	15'h52a: q<=8'h11;
	15'h52b: q<=8'h20;
	15'h52c: q<=8'h05;
	15'h52d: q<=8'h03;
	15'h52e: q<=8'h02;
	15'h52f: q<=8'h02;
	15'h530: q<=8'h02;
	15'h531: q<=8'h02;
	15'h532: q<=8'h02;
	15'h533: q<=8'h02;
	15'h534: q<=8'h02;
	15'h535: q<=8'h02;
	15'h536: q<=8'h02;
	15'h537: q<=8'h02;
	15'h538: q<=8'h02;
	15'h539: q<=8'h03;
	15'h53a: q<=8'h04;
	15'h53b: q<=8'h02;
	15'h53c: q<=8'h02;
	15'h53d: q<=8'h21;
	15'h53e: q<=8'h63;
	15'h53f: q<=8'h03;
	15'h540: q<=8'h00;
	15'h541: q<=8'h02;
	15'h542: q<=8'h0b;
	15'h543: q<=8'h10;
	15'h544: q<=8'h01;
	15'h545: q<=8'h02;
	15'h546: q<=8'h16;
	15'h547: q<=8'h19;
	15'h548: q<=8'h01;
	15'h549: q<=8'h02;
	15'h54a: q<=8'h1b;
	15'h54b: q<=8'h63;
	15'h54c: q<=8'h01;
	15'h54d: q<=8'h00;
	15'h54e: q<=8'h02;
	15'h54f: q<=8'h0b;
	15'h550: q<=8'h10;
	15'h551: q<=8'h01;
	15'h552: q<=8'h02;
	15'h553: q<=8'h16;
	15'h554: q<=8'h19;
	15'h555: q<=8'h01;
	15'h556: q<=8'h02;
	15'h557: q<=8'h1b;
	15'h558: q<=8'h20;
	15'h559: q<=8'h01;
	15'h55a: q<=8'h02;
	15'h55b: q<=8'h21;
	15'h55c: q<=8'h27;
	15'h55d: q<=8'h04;
	15'h55e: q<=8'h02;
	15'h55f: q<=8'h28;
	15'h560: q<=8'h63;
	15'h561: q<=8'h03;
	15'h562: q<=8'h00;
	15'h563: q<=8'h04;
	15'h564: q<=8'h11;
	15'h565: q<=8'h12;
	15'h566: q<=8'h28;
	15'h567: q<=8'h14;
	15'h568: q<=8'h0c;
	15'h569: q<=8'h13;
	15'h56a: q<=8'h20;
	15'h56b: q<=8'h14;
	15'h56c: q<=8'h28;
	15'h56d: q<=8'h08;
	15'h56e: q<=8'h21;
	15'h56f: q<=8'h27;
	15'h570: q<=8'h14;
	15'h571: q<=8'hff;
	15'h572: q<=8'h0c;
	15'h573: q<=8'h28;
	15'h574: q<=8'h63;
	15'h575: q<=8'h14;
	15'h576: q<=8'h0a;
	15'h577: q<=8'h00;
	15'h578: q<=8'h0c;
	15'h579: q<=8'h11;
	15'h57a: q<=8'h20;
	15'h57b: q<=8'h00;
	15'h57c: q<=8'h40;
	15'h57d: q<=8'h0c;
	15'h57e: q<=8'h21;
	15'h57f: q<=8'h30;
	15'h580: q<=8'h40;
	15'h581: q<=8'hc0;
	15'h582: q<=8'h02;
	15'h583: q<=8'h31;
	15'h584: q<=8'h63;
	15'h585: q<=8'hc0;
	15'h586: q<=8'h00;
	15'h587: q<=8'h02;
	15'h588: q<=8'h01;
	15'h589: q<=8'h10;
	15'h58a: q<=8'hdc;
	15'h58b: q<=8'h02;
	15'h58c: q<=8'h11;
	15'h58d: q<=8'h27;
	15'h58e: q<=8'hc0;
	15'h58f: q<=8'h08;
	15'h590: q<=8'h28;
	15'h591: q<=8'h40;
	15'h592: q<=8'hc0;
	15'h593: q<=8'h01;
	15'h594: q<=8'h02;
	15'h595: q<=8'h41;
	15'h596: q<=8'h63;
	15'h597: q<=8'he6;
	15'h598: q<=8'h02;
	15'h599: q<=8'h01;
	15'h59a: q<=8'h63;
	15'h59b: q<=8'h06;
	15'h59c: q<=8'h06;
	15'h59d: q<=8'h01;
	15'h59e: q<=8'h63;
	15'h59f: q<=8'h00;
	15'h5a0: q<=8'h00;
	15'h5a1: q<=8'h00;
	15'h5a2: q<=8'he0;
	15'h5a3: q<=8'hd8;
	15'h5a4: q<=8'hd4;
	15'h5a5: q<=8'hd0;
	15'h5a6: q<=8'hc8;
	15'h5a7: q<=8'hc0;
	15'h5a8: q<=8'hb8;
	15'h5a9: q<=8'hb0;
	15'h5aa: q<=8'ha8;
	15'h5ab: q<=8'ha0;
	15'h5ac: q<=8'ha0;
	15'h5ad: q<=8'ha0;
	15'h5ae: q<=8'ha8;
	15'h5af: q<=8'ha0;
	15'h5b0: q<=8'h9c;
	15'h5b1: q<=8'h9a;
	15'h5b2: q<=8'h98;
	15'h5b3: q<=8'h04;
	15'h5b4: q<=8'h01;
	15'h5b5: q<=8'h10;
	15'h5b6: q<=8'h0a;
	15'h5b7: q<=8'h0c;
	15'h5b8: q<=8'h0f;
	15'h5b9: q<=8'h11;
	15'h5ba: q<=8'h14;
	15'h5bb: q<=8'h16;
	15'h5bc: q<=8'h14;
	15'h5bd: q<=8'h18;
	15'h5be: q<=8'h1b;
	15'h5bf: q<=8'h1d;
	15'h5c0: q<=8'h1b;
	15'h5c1: q<=8'h18;
	15'h5c2: q<=8'h1a;
	15'h5c3: q<=8'h1c;
	15'h5c4: q<=8'h1e;
	15'h5c5: q<=8'h1b;
	15'h5c6: q<=8'h08;
	15'h5c7: q<=8'h11;
	15'h5c8: q<=8'h1a;
	15'h5c9: q<=8'h14;
	15'h5ca: q<=8'h01;
	15'h5cb: q<=8'h02;
	15'h5cc: q<=8'h1b;
	15'h5cd: q<=8'h27;
	15'h5ce: q<=8'h1b;
	15'h5cf: q<=8'h08;
	15'h5d0: q<=8'h28;
	15'h5d1: q<=8'h30;
	15'h5d2: q<=8'h1d;
	15'h5d3: q<=8'h01;
	15'h5d4: q<=8'h08;
	15'h5d5: q<=8'h31;
	15'h5d6: q<=8'h40;
	15'h5d7: q<=8'h1f;
	15'h5d8: q<=8'h01;
	15'h5d9: q<=8'h08;
	15'h5da: q<=8'h41;
	15'h5db: q<=8'h50;
	15'h5dc: q<=8'h23;
	15'h5dd: q<=8'h01;
	15'h5de: q<=8'h08;
	15'h5df: q<=8'h51;
	15'h5e0: q<=8'h63;
	15'h5e1: q<=8'h2b;
	15'h5e2: q<=8'h01;
	15'h5e3: q<=8'h02;
	15'h5e4: q<=8'h01;
	15'h5e5: q<=8'h14;
	15'h5e6: q<=8'h02;
	15'h5e7: q<=8'h02;
	15'h5e8: q<=8'h15;
	15'h5e9: q<=8'h20;
	15'h5ea: q<=8'h02;
	15'h5eb: q<=8'h02;
	15'h5ec: q<=8'h21;
	15'h5ed: q<=8'h63;
	15'h5ee: q<=8'h03;
	15'h5ef: q<=8'h02;
	15'h5f0: q<=8'h3c;
	15'h5f1: q<=8'h63;
	15'h5f2: q<=8'h40;
	15'h5f3: q<=8'h00;
	15'h5f4: q<=8'h06;
	15'h5f5: q<=8'h01;
	15'h5f6: q<=8'h63;
	15'h5f7: q<=8'h07;
	15'h5f8: q<=8'h0b;
	15'h5f9: q<=8'h19;
	15'h5fa: q<=8'h24;
	15'h5fb: q<=8'h53;
	15'h5fc: q<=8'h0b;
	15'h5fd: q<=8'h24;
	15'h5fe: q<=8'h19;
	15'h5ff: q<=8'h53;
	15'h600: q<=8'h87;
	15'h601: q<=8'h24;
	15'h602: q<=8'h19;
	15'h603: q<=8'h53;
	15'h604: q<=8'h07;
	15'h605: q<=8'h87;
	15'h606: q<=8'h24;
	15'h607: q<=8'hef;
	15'h608: q<=8'h95;
	15'h609: q<=8'h6d;
	15'h60a: q<=8'h01;
	15'h60b: q<=8'he3;
	15'h60c: q<=8'h95;
	15'h60d: q<=8'hb3;
	15'h60e: q<=8'h00;
	15'h60f: q<=8'hfa;
	15'h610: q<=8'h93;
	15'h611: q<=8'h19;
	15'h612: q<=8'h01;
	15'h613: q<=8'h07;
	15'h614: q<=8'h94;
	15'h615: q<=8'h1a;
	15'h616: q<=8'h01;
	15'h617: q<=8'hcd;
	15'h618: q<=8'h94;
	15'h619: q<=8'h29;
	15'h61a: q<=8'h01;
	15'h61b: q<=8'hd6;
	15'h61c: q<=8'h94;
	15'h61d: q<=8'h2e;
	15'h61e: q<=8'h01;
	15'h61f: q<=8'h20;
	15'h620: q<=8'h95;
	15'h621: q<=8'h2a;
	15'h622: q<=8'h01;
	15'h623: q<=8'h29;
	15'h624: q<=8'h95;
	15'h625: q<=8'h2f;
	15'h626: q<=8'h01;
	15'h627: q<=8'heb;
	15'h628: q<=8'h94;
	15'h629: q<=8'h2b;
	15'h62a: q<=8'h01;
	15'h62b: q<=8'h03;
	15'h62c: q<=8'h95;
	15'h62d: q<=8'h30;
	15'h62e: q<=8'h01;
	15'h62f: q<=8'h89;
	15'h630: q<=8'h94;
	15'h631: q<=8'h2c;
	15'h632: q<=8'h01;
	15'h633: q<=8'ha5;
	15'h634: q<=8'h94;
	15'h635: q<=8'h31;
	15'h636: q<=8'h01;
	15'h637: q<=8'h41;
	15'h638: q<=8'h95;
	15'h639: q<=8'h2d;
	15'h63a: q<=8'h01;
	15'h63b: q<=8'h4e;
	15'h63c: q<=8'h95;
	15'h63d: q<=8'h32;
	15'h63e: q<=8'h01;
	15'h63f: q<=8'h5d;
	15'h640: q<=8'h94;
	15'h641: q<=8'h57;
	15'h642: q<=8'h01;
	15'h643: q<=8'h69;
	15'h644: q<=8'h94;
	15'h645: q<=8'h47;
	15'h646: q<=8'h01;
	15'h647: q<=8'h75;
	15'h648: q<=8'h94;
	15'h649: q<=8'h4b;
	15'h64a: q<=8'h01;
	15'h64b: q<=8'h81;
	15'h64c: q<=8'h94;
	15'h64d: q<=8'h4c;
	15'h64e: q<=8'h01;
	15'h64f: q<=8'h98;
	15'h650: q<=8'h95;
	15'h651: q<=8'h1c;
	15'h652: q<=8'h01;
	15'h653: q<=8'hb3;
	15'h654: q<=8'h95;
	15'h655: q<=8'h5b;
	15'h656: q<=8'h01;
	15'h657: q<=8'h9c;
	15'h658: q<=8'h95;
	15'h659: q<=8'h5a;
	15'h65a: q<=8'h01;
	15'h65b: q<=8'h63;
	15'h65c: q<=8'h95;
	15'h65d: q<=8'hb2;
	15'h65e: q<=8'h00;
	15'h65f: q<=8'hf4;
	15'h660: q<=8'h95;
	15'h661: q<=8'h5d;
	15'h662: q<=8'h01;
	15'h663: q<=8'h4d;
	15'h664: q<=8'h94;
	15'h665: q<=8'h63;
	15'h666: q<=8'h01;
	15'h667: q<=8'h49;
	15'h668: q<=8'h94;
	15'h669: q<=8'h20;
	15'h66a: q<=8'h01;
	15'h66b: q<=8'h1b;
	15'h66c: q<=8'h94;
	15'h66d: q<=8'h60;
	15'h66e: q<=8'h01;
	15'h66f: q<=8'h78;
	15'h670: q<=8'h95;
	15'h671: q<=8'h59;
	15'h672: q<=8'h01;
	15'h673: q<=8'h87;
	15'h674: q<=8'h95;
	15'h675: q<=8'h5f;
	15'h676: q<=8'h01;
	15'h677: q<=8'hae;
	15'h678: q<=8'h5e;
	15'h679: q<=8'h01;
	15'h67a: q<=8'hbd;
	15'h67b: q<=8'h90;
	15'h67c: q<=8'h96;
	15'h67d: q<=8'h48;
	15'h67e: q<=8'hbd;
	15'h67f: q<=8'h8f;
	15'h680: q<=8'h96;
	15'h681: q<=8'h48;
	15'h682: q<=8'h60;
	15'h683: q<=8'hae;
	15'h684: q<=8'h5e;
	15'h685: q<=8'h01;
	15'h686: q<=8'hbd;
	15'h687: q<=8'h9e;
	15'h688: q<=8'h96;
	15'h689: q<=8'h48;
	15'h68a: q<=8'hbd;
	15'h68b: q<=8'h9d;
	15'h68c: q<=8'h96;
	15'h68d: q<=8'h48;
	15'h68e: q<=8'h60;
	15'h68f: q<=8'h00;
	15'h690: q<=8'h00;
	15'h691: q<=8'hc3;
	15'h692: q<=8'h96;
	15'h693: q<=8'hb6;
	15'h694: q<=8'h96;
	15'h695: q<=8'haa;
	15'h696: q<=8'h96;
	15'h697: q<=8'he1;
	15'h698: q<=8'h96;
	15'h699: q<=8'hda;
	15'h69a: q<=8'h96;
	15'h69b: q<=8'hff;
	15'h69c: q<=8'h96;
	15'h69d: q<=8'h00;
	15'h69e: q<=8'h00;
	15'h69f: q<=8'hc7;
	15'h6a0: q<=8'h96;
	15'h6a1: q<=8'hca;
	15'h6a2: q<=8'h96;
	15'h6a3: q<=8'hca;
	15'h6a4: q<=8'h96;
	15'h6a5: q<=8'hc6;
	15'h6a6: q<=8'h96;
	15'h6a7: q<=8'hc7;
	15'h6a8: q<=8'h96;
	15'h6a9: q<=8'hc6;
	15'h6aa: q<=8'h96;
	15'h6ab: q<=8'ha5;
	15'h6ac: q<=8'h2b;
	15'h6ad: q<=8'h38;
	15'h6ae: q<=8'he9;
	15'h6af: q<=8'h01;
	15'h6b0: q<=8'h29;
	15'h6b1: q<=8'h0f;
	15'h6b2: q<=8'h18;
	15'h6b3: q<=8'h69;
	15'h6b4: q<=8'h01;
	15'h6b5: q<=8'h10;
	15'h6b6: q<=8'h02;
	15'h6b7: q<=8'ha5;
	15'h6b8: q<=8'h2b;
	15'h6b9: q<=8'h84;
	15'h6ba: q<=8'h29;
	15'h6bb: q<=8'h88;
	15'h6bc: q<=8'h88;
	15'h6bd: q<=8'h38;
	15'h6be: q<=8'hf1;
	15'h6bf: q<=8'h2c;
	15'h6c0: q<=8'h18;
	15'h6c1: q<=8'h65;
	15'h6c2: q<=8'h29;
	15'h6c3: q<=8'ha8;
	15'h6c4: q<=8'hb1;
	15'h6c5: q<=8'h2c;
	15'h6c6: q<=8'h60;
	15'h6c7: q<=8'hc8;
	15'h6c8: q<=8'hc8;
	15'h6c9: q<=8'hc8;
	15'h6ca: q<=8'h60;
	15'h6cb: q<=8'hb1;
	15'h6cc: q<=8'h2c;
	15'h6cd: q<=8'h88;
	15'h6ce: q<=8'h38;
	15'h6cf: q<=8'hf1;
	15'h6d0: q<=8'h2c;
	15'h6d1: q<=8'h85;
	15'h6d2: q<=8'h29;
	15'h6d3: q<=8'h98;
	15'h6d4: q<=8'h38;
	15'h6d5: q<=8'h65;
	15'h6d6: q<=8'h29;
	15'h6d7: q<=8'ha8;
	15'h6d8: q<=8'hc8;
	15'h6d9: q<=8'hc8;
	15'h6da: q<=8'h60;
	15'h6db: q<=8'hb1;
	15'h6dc: q<=8'h2c;
	15'h6dd: q<=8'h18;
	15'h6de: q<=8'h6d;
	15'h6df: q<=8'h60;
	15'h6e0: q<=8'h01;
	15'h6e1: q<=8'h60;
	15'h6e2: q<=8'h20;
	15'h6e3: q<=8'hf4;
	15'h6e4: q<=8'h96;
	15'h6e5: q<=8'haa;
	15'h6e6: q<=8'hb1;
	15'h6e7: q<=8'h2c;
	15'h6e8: q<=8'hc8;
	15'h6e9: q<=8'he0;
	15'h6ea: q<=8'h00;
	15'h6eb: q<=8'hf0;
	15'h6ec: q<=8'h06;
	15'h6ed: q<=8'h18;
	15'h6ee: q<=8'h71;
	15'h6ef: q<=8'h2c;
	15'h6f0: q<=8'hca;
	15'h6f1: q<=8'hd0;
	15'h6f2: q<=8'hfa;
	15'h6f3: q<=8'h60;
	15'h6f4: q<=8'ha5;
	15'h6f5: q<=8'h2b;
	15'h6f6: q<=8'h84;
	15'h6f7: q<=8'h29;
	15'h6f8: q<=8'h88;
	15'h6f9: q<=8'h88;
	15'h6fa: q<=8'h38;
	15'h6fb: q<=8'hf1;
	15'h6fc: q<=8'h2c;
	15'h6fd: q<=8'hc8;
	15'h6fe: q<=8'hc8;
	15'h6ff: q<=8'h60;
	15'h700: q<=8'h20;
	15'h701: q<=8'hf4;
	15'h702: q<=8'h96;
	15'h703: q<=8'h29;
	15'h704: q<=8'h01;
	15'h705: q<=8'hf0;
	15'h706: q<=8'h01;
	15'h707: q<=8'hc8;
	15'h708: q<=8'hb1;
	15'h709: q<=8'h2c;
	15'h70a: q<=8'h60;
	15'h70b: q<=8'h20;
	15'h70c: q<=8'h49;
	15'h70d: q<=8'h97;
	15'h70e: q<=8'h20;
	15'h70f: q<=8'h3f;
	15'h710: q<=8'ha2;
	15'h711: q<=8'h20;
	15'h712: q<=8'h3a;
	15'h713: q<=8'ha8;
	15'h714: q<=8'h20;
	15'h715: q<=8'ha2;
	15'h716: q<=8'h98;
	15'h717: q<=8'h20;
	15'h718: q<=8'h1e;
	15'h719: q<=8'h9b;
	15'h71a: q<=8'h20;
	15'h71b: q<=8'h8f;
	15'h71c: q<=8'ha1;
	15'h71d: q<=8'h20;
	15'h71e: q<=8'ha6;
	15'h71f: q<=8'ha2;
	15'h720: q<=8'h20;
	15'h721: q<=8'h54;
	15'h722: q<=8'ha4;
	15'h723: q<=8'h20;
	15'h724: q<=8'h16;
	15'h725: q<=8'ha4;
	15'h726: q<=8'h4c;
	15'h727: q<=8'h04;
	15'h728: q<=8'ha5;
	15'h729: q<=8'had;
	15'h72a: q<=8'h23;
	15'h72b: q<=8'h01;
	15'h72c: q<=8'h29;
	15'h72d: q<=8'h7f;
	15'h72e: q<=8'h8d;
	15'h72f: q<=8'h23;
	15'h730: q<=8'h01;
	15'h731: q<=8'h20;
	15'h732: q<=8'h49;
	15'h733: q<=8'h97;
	15'h734: q<=8'h20;
	15'h735: q<=8'hf8;
	15'h736: q<=8'h97;
	15'h737: q<=8'h20;
	15'h738: q<=8'h16;
	15'h739: q<=8'ha4;
	15'h73a: q<=8'h20;
	15'h73b: q<=8'h3f;
	15'h73c: q<=8'ha2;
	15'h73d: q<=8'h20;
	15'h73e: q<=8'h8f;
	15'h73f: q<=8'ha1;
	15'h740: q<=8'had;
	15'h741: q<=8'h01;
	15'h742: q<=8'h02;
	15'h743: q<=8'h10;
	15'h744: q<=8'h03;
	15'h745: q<=8'h20;
	15'h746: q<=8'h04;
	15'h747: q<=8'ha5;
	15'h748: q<=8'h60;
	15'h749: q<=8'had;
	15'h74a: q<=8'h01;
	15'h74b: q<=8'h02;
	15'h74c: q<=8'h10;
	15'h74d: q<=8'h01;
	15'h74e: q<=8'h60;
	15'h74f: q<=8'ha2;
	15'h750: q<=8'h00;
	15'h751: q<=8'ha5;
	15'h752: q<=8'h05;
	15'h753: q<=8'h30;
	15'h754: q<=8'h06;
	15'h755: q<=8'h20;
	15'h756: q<=8'hc5;
	15'h757: q<=8'h97;
	15'h758: q<=8'hb8;
	15'h759: q<=8'h50;
	15'h75a: q<=8'h15;
	15'h75b: q<=8'ha5;
	15'h75c: q<=8'h50;
	15'h75d: q<=8'h10;
	15'h75e: q<=8'h09;
	15'h75f: q<=8'hc9;
	15'h760: q<=8'he1;
	15'h761: q<=8'hb0;
	15'h762: q<=8'h02;
	15'h763: q<=8'ha9;
	15'h764: q<=8'he1;
	15'h765: q<=8'hb8;
	15'h766: q<=8'h50;
	15'h767: q<=8'h06;
	15'h768: q<=8'hc9;
	15'h769: q<=8'h1f;
	15'h76a: q<=8'h90;
	15'h76b: q<=8'h02;
	15'h76c: q<=8'ha9;
	15'h76d: q<=8'h1f;
	15'h76e: q<=8'h86;
	15'h76f: q<=8'h50;
	15'h770: q<=8'h85;
	15'h771: q<=8'h2b;
	15'h772: q<=8'h49;
	15'h773: q<=8'hff;
	15'h774: q<=8'h38;
	15'h775: q<=8'h65;
	15'h776: q<=8'h51;
	15'h777: q<=8'h85;
	15'h778: q<=8'h2c;
	15'h779: q<=8'hae;
	15'h77a: q<=8'h11;
	15'h77b: q<=8'h01;
	15'h77c: q<=8'hf0;
	15'h77d: q<=8'h1f;
	15'h77e: q<=8'hc9;
	15'h77f: q<=8'hf0;
	15'h780: q<=8'h90;
	15'h781: q<=8'h04;
	15'h782: q<=8'ha9;
	15'h783: q<=8'hef;
	15'h784: q<=8'h85;
	15'h785: q<=8'h2c;
	15'h786: q<=8'h45;
	15'h787: q<=8'h2b;
	15'h788: q<=8'h10;
	15'h789: q<=8'h13;
	15'h78a: q<=8'ha5;
	15'h78b: q<=8'h2c;
	15'h78c: q<=8'h45;
	15'h78d: q<=8'h51;
	15'h78e: q<=8'h10;
	15'h78f: q<=8'h0d;
	15'h790: q<=8'ha5;
	15'h791: q<=8'h51;
	15'h792: q<=8'h30;
	15'h793: q<=8'h05;
	15'h794: q<=8'ha9;
	15'h795: q<=8'h00;
	15'h796: q<=8'hb8;
	15'h797: q<=8'h50;
	15'h798: q<=8'h02;
	15'h799: q<=8'ha9;
	15'h79a: q<=8'hef;
	15'h79b: q<=8'h85;
	15'h79c: q<=8'h2c;
	15'h79d: q<=8'ha5;
	15'h79e: q<=8'h2c;
	15'h79f: q<=8'h4a;
	15'h7a0: q<=8'h4a;
	15'h7a1: q<=8'h4a;
	15'h7a2: q<=8'h4a;
	15'h7a3: q<=8'h85;
	15'h7a4: q<=8'h2a;
	15'h7a5: q<=8'h18;
	15'h7a6: q<=8'h69;
	15'h7a7: q<=8'h01;
	15'h7a8: q<=8'h29;
	15'h7a9: q<=8'h0f;
	15'h7aa: q<=8'h85;
	15'h7ab: q<=8'h2b;
	15'h7ac: q<=8'ha5;
	15'h7ad: q<=8'h2a;
	15'h7ae: q<=8'hcd;
	15'h7af: q<=8'h00;
	15'h7b0: q<=8'h02;
	15'h7b1: q<=8'hf0;
	15'h7b2: q<=8'h03;
	15'h7b3: q<=8'h20;
	15'h7b4: q<=8'hb5;
	15'h7b5: q<=8'hcc;
	15'h7b6: q<=8'ha5;
	15'h7b7: q<=8'h2a;
	15'h7b8: q<=8'h8d;
	15'h7b9: q<=8'h00;
	15'h7ba: q<=8'h02;
	15'h7bb: q<=8'ha5;
	15'h7bc: q<=8'h2b;
	15'h7bd: q<=8'h8d;
	15'h7be: q<=8'h01;
	15'h7bf: q<=8'h02;
	15'h7c0: q<=8'ha5;
	15'h7c1: q<=8'h2c;
	15'h7c2: q<=8'h85;
	15'h7c3: q<=8'h51;
	15'h7c4: q<=8'h60;
	15'h7c5: q<=8'ha9;
	15'h7c6: q<=8'hff;
	15'h7c7: q<=8'h85;
	15'h7c8: q<=8'h29;
	15'h7c9: q<=8'h85;
	15'h7ca: q<=8'h2a;
	15'h7cb: q<=8'hae;
	15'h7cc: q<=8'h1c;
	15'h7cd: q<=8'h01;
	15'h7ce: q<=8'hbd;
	15'h7cf: q<=8'hdf;
	15'h7d0: q<=8'h02;
	15'h7d1: q<=8'hf0;
	15'h7d2: q<=8'h08;
	15'h7d3: q<=8'hc5;
	15'h7d4: q<=8'h29;
	15'h7d5: q<=8'hb0;
	15'h7d6: q<=8'h04;
	15'h7d7: q<=8'h85;
	15'h7d8: q<=8'h29;
	15'h7d9: q<=8'h86;
	15'h7da: q<=8'h2a;
	15'h7db: q<=8'hca;
	15'h7dc: q<=8'h10;
	15'h7dd: q<=8'hf0;
	15'h7de: q<=8'ha6;
	15'h7df: q<=8'h2a;
	15'h7e0: q<=8'h30;
	15'h7e1: q<=8'h15;
	15'h7e2: q<=8'hbd;
	15'h7e3: q<=8'hb9;
	15'h7e4: q<=8'h02;
	15'h7e5: q<=8'hac;
	15'h7e6: q<=8'h00;
	15'h7e7: q<=8'h02;
	15'h7e8: q<=8'h20;
	15'h7e9: q<=8'ha6;
	15'h7ea: q<=8'ha7;
	15'h7eb: q<=8'ha8;
	15'h7ec: q<=8'hf0;
	15'h7ed: q<=8'h09;
	15'h7ee: q<=8'h30;
	15'h7ef: q<=8'h05;
	15'h7f0: q<=8'ha9;
	15'h7f1: q<=8'hf7;
	15'h7f2: q<=8'hb8;
	15'h7f3: q<=8'h50;
	15'h7f4: q<=8'h02;
	15'h7f5: q<=8'ha9;
	15'h7f6: q<=8'h09;
	15'h7f7: q<=8'h60;
	15'h7f8: q<=8'had;
	15'h7f9: q<=8'h01;
	15'h7fa: q<=8'h02;
	15'h7fb: q<=8'h10;
	15'h7fc: q<=8'h01;
	15'h7fd: q<=8'h60;
	15'h7fe: q<=8'had;
	15'h7ff: q<=8'h06;
	15'h800: q<=8'h01;
	15'h801: q<=8'h30;
	15'h802: q<=8'h01;
	15'h803: q<=8'h60;
	15'h804: q<=8'had;
	15'h805: q<=8'h02;
	15'h806: q<=8'h02;
	15'h807: q<=8'hc9;
	15'h808: q<=8'h10;
	15'h809: q<=8'hd0;
	15'h80a: q<=8'h03;
	15'h80b: q<=8'h20;
	15'h80c: q<=8'hee;
	15'h80d: q<=8'hcc;
	15'h80e: q<=8'had;
	15'h80f: q<=8'h07;
	15'h810: q<=8'h01;
	15'h811: q<=8'h18;
	15'h812: q<=8'h6d;
	15'h813: q<=8'h04;
	15'h814: q<=8'h01;
	15'h815: q<=8'h8d;
	15'h816: q<=8'h07;
	15'h817: q<=8'h01;
	15'h818: q<=8'had;
	15'h819: q<=8'h02;
	15'h81a: q<=8'h02;
	15'h81b: q<=8'h6d;
	15'h81c: q<=8'h05;
	15'h81d: q<=8'h01;
	15'h81e: q<=8'h8d;
	15'h81f: q<=8'h02;
	15'h820: q<=8'h02;
	15'h821: q<=8'hb0;
	15'h822: q<=8'h02;
	15'h823: q<=8'hc9;
	15'h824: q<=8'hf0;
	15'h825: q<=8'h90;
	15'h826: q<=8'h0c;
	15'h827: q<=8'ha9;
	15'h828: q<=8'h0e;
	15'h829: q<=8'h85;
	15'h82a: q<=8'h00;
	15'h82b: q<=8'h20;
	15'h82c: q<=8'hf2;
	15'h82d: q<=8'hcc;
	15'h82e: q<=8'ha9;
	15'h82f: q<=8'hff;
	15'h830: q<=8'h8d;
	15'h831: q<=8'h02;
	15'h832: q<=8'h02;
	15'h833: q<=8'had;
	15'h834: q<=8'h02;
	15'h835: q<=8'h02;
	15'h836: q<=8'hc9;
	15'h837: q<=8'h50;
	15'h838: q<=8'h90;
	15'h839: q<=8'h08;
	15'h83a: q<=8'had;
	15'h83b: q<=8'h15;
	15'h83c: q<=8'h01;
	15'h83d: q<=8'hd0;
	15'h83e: q<=8'h03;
	15'h83f: q<=8'h20;
	15'h840: q<=8'hbd;
	15'h841: q<=8'ha7;
	15'h842: q<=8'ha5;
	15'h843: q<=8'h5c;
	15'h844: q<=8'h18;
	15'h845: q<=8'h6d;
	15'h846: q<=8'h04;
	15'h847: q<=8'h01;
	15'h848: q<=8'h85;
	15'h849: q<=8'h5c;
	15'h84a: q<=8'ha5;
	15'h84b: q<=8'h5f;
	15'h84c: q<=8'h6d;
	15'h84d: q<=8'h05;
	15'h84e: q<=8'h01;
	15'h84f: q<=8'h90;
	15'h850: q<=8'h02;
	15'h851: q<=8'he6;
	15'h852: q<=8'h5b;
	15'h853: q<=8'hc5;
	15'h854: q<=8'h5f;
	15'h855: q<=8'hf0;
	15'h856: q<=8'h03;
	15'h857: q<=8'hee;
	15'h858: q<=8'h14;
	15'h859: q<=8'h01;
	15'h85a: q<=8'h85;
	15'h85b: q<=8'h5f;
	15'h85c: q<=8'ha5;
	15'h85d: q<=8'h9f;
	15'h85e: q<=8'h0a;
	15'h85f: q<=8'h0a;
	15'h860: q<=8'hc9;
	15'h861: q<=8'h30;
	15'h862: q<=8'h90;
	15'h863: q<=8'h02;
	15'h864: q<=8'ha9;
	15'h865: q<=8'h30;
	15'h866: q<=8'h18;
	15'h867: q<=8'h69;
	15'h868: q<=8'h20;
	15'h869: q<=8'h18;
	15'h86a: q<=8'h6d;
	15'h86b: q<=8'h04;
	15'h86c: q<=8'h01;
	15'h86d: q<=8'h8d;
	15'h86e: q<=8'h04;
	15'h86f: q<=8'h01;
	15'h870: q<=8'had;
	15'h871: q<=8'h05;
	15'h872: q<=8'h01;
	15'h873: q<=8'h69;
	15'h874: q<=8'h00;
	15'h875: q<=8'h8d;
	15'h876: q<=8'h05;
	15'h877: q<=8'h01;
	15'h878: q<=8'had;
	15'h879: q<=8'h02;
	15'h87a: q<=8'h02;
	15'h87b: q<=8'hc9;
	15'h87c: q<=8'hf0;
	15'h87d: q<=8'hb0;
	15'h87e: q<=8'h22;
	15'h87f: q<=8'ha2;
	15'h880: q<=8'h0f;
	15'h881: q<=8'hbd;
	15'h882: q<=8'hac;
	15'h883: q<=8'h03;
	15'h884: q<=8'hf0;
	15'h885: q<=8'h18;
	15'h886: q<=8'hec;
	15'h887: q<=8'h00;
	15'h888: q<=8'h02;
	15'h889: q<=8'hd0;
	15'h88a: q<=8'h13;
	15'h88b: q<=8'hcd;
	15'h88c: q<=8'h02;
	15'h88d: q<=8'h02;
	15'h88e: q<=8'hb0;
	15'h88f: q<=8'h0e;
	15'h890: q<=8'h20;
	15'h891: q<=8'h06;
	15'h892: q<=8'hcd;
	15'h893: q<=8'h20;
	15'h894: q<=8'h47;
	15'h895: q<=8'ha3;
	15'h896: q<=8'ha9;
	15'h897: q<=8'h00;
	15'h898: q<=8'h8d;
	15'h899: q<=8'h15;
	15'h89a: q<=8'h01;
	15'h89b: q<=8'h20;
	15'h89c: q<=8'h8f;
	15'h89d: q<=8'h92;
	15'h89e: q<=8'hca;
	15'h89f: q<=8'h10;
	15'h8a0: q<=8'he0;
	15'h8a1: q<=8'h60;
	15'h8a2: q<=8'ha0;
	15'h8a3: q<=8'h00;
	15'h8a4: q<=8'h8c;
	15'h8a5: q<=8'h4f;
	15'h8a6: q<=8'h01;
	15'h8a7: q<=8'had;
	15'h8a8: q<=8'h08;
	15'h8a9: q<=8'h01;
	15'h8aa: q<=8'h18;
	15'h8ab: q<=8'h6d;
	15'h8ac: q<=8'h09;
	15'h8ad: q<=8'h01;
	15'h8ae: q<=8'hcd;
	15'h8af: q<=8'h1c;
	15'h8b0: q<=8'h01;
	15'h8b1: q<=8'h90;
	15'h8b2: q<=8'h04;
	15'h8b3: q<=8'hf0;
	15'h8b4: q<=8'h02;
	15'h8b5: q<=8'ha0;
	15'h8b6: q<=8'hff;
	15'h8b7: q<=8'had;
	15'h8b8: q<=8'h25;
	15'h8b9: q<=8'h01;
	15'h8ba: q<=8'hf0;
	15'h8bb: q<=8'h02;
	15'h8bc: q<=8'ha0;
	15'h8bd: q<=8'hff;
	15'h8be: q<=8'h84;
	15'h8bf: q<=8'h2f;
	15'h8c0: q<=8'ha2;
	15'h8c1: q<=8'h3f;
	15'h8c2: q<=8'hbd;
	15'h8c3: q<=8'h43;
	15'h8c4: q<=8'h02;
	15'h8c5: q<=8'hf0;
	15'h8c6: q<=8'h52;
	15'h8c7: q<=8'h24;
	15'h8c8: q<=8'h2f;
	15'h8c9: q<=8'h30;
	15'h8ca: q<=8'h23;
	15'h8cb: q<=8'h38;
	15'h8cc: q<=8'he9;
	15'h8cd: q<=8'h01;
	15'h8ce: q<=8'h9d;
	15'h8cf: q<=8'h43;
	15'h8d0: q<=8'h02;
	15'h8d1: q<=8'hd0;
	15'h8d2: q<=8'h06;
	15'h8d3: q<=8'h20;
	15'h8d4: q<=8'h23;
	15'h8d5: q<=8'h99;
	15'h8d6: q<=8'hb8;
	15'h8d7: q<=8'h50;
	15'h8d8: q<=8'h15;
	15'h8d9: q<=8'hc9;
	15'h8da: q<=8'h3f;
	15'h8db: q<=8'hd0;
	15'h8dc: q<=8'h11;
	15'h8dd: q<=8'hbc;
	15'h8de: q<=8'h03;
	15'h8df: q<=8'h02;
	15'h8e0: q<=8'had;
	15'h8e1: q<=8'h4f;
	15'h8e2: q<=8'h01;
	15'h8e3: q<=8'h0d;
	15'h8e4: q<=8'h4f;
	15'h8e5: q<=8'h01;
	15'h8e6: q<=8'h39;
	15'h8e7: q<=8'h38;
	15'h8e8: q<=8'hca;
	15'h8e9: q<=8'hf0;
	15'h8ea: q<=8'h03;
	15'h8eb: q<=8'hfe;
	15'h8ec: q<=8'h43;
	15'h8ed: q<=8'h02;
	15'h8ee: q<=8'hbd;
	15'h8ef: q<=8'h43;
	15'h8f0: q<=8'h02;
	15'h8f1: q<=8'hc9;
	15'h8f2: q<=8'h40;
	15'h8f3: q<=8'h90;
	15'h8f4: q<=8'h14;
	15'h8f5: q<=8'ha5;
	15'h8f6: q<=8'h03;
	15'h8f7: q<=8'h29;
	15'h8f8: q<=8'h01;
	15'h8f9: q<=8'hd0;
	15'h8fa: q<=8'h0b;
	15'h8fb: q<=8'hbd;
	15'h8fc: q<=8'h03;
	15'h8fd: q<=8'h02;
	15'h8fe: q<=8'h18;
	15'h8ff: q<=8'h69;
	15'h900: q<=8'h01;
	15'h901: q<=8'h29;
	15'h902: q<=8'h0f;
	15'h903: q<=8'h9d;
	15'h904: q<=8'h03;
	15'h905: q<=8'h02;
	15'h906: q<=8'hb8;
	15'h907: q<=8'h50;
	15'h908: q<=8'h10;
	15'h909: q<=8'hc9;
	15'h90a: q<=8'h20;
	15'h90b: q<=8'h90;
	15'h90c: q<=8'h0c;
	15'h90d: q<=8'hbc;
	15'h90e: q<=8'h03;
	15'h90f: q<=8'h02;
	15'h910: q<=8'hb9;
	15'h911: q<=8'h38;
	15'h912: q<=8'hca;
	15'h913: q<=8'h0d;
	15'h914: q<=8'h4f;
	15'h915: q<=8'h01;
	15'h916: q<=8'h8d;
	15'h917: q<=8'h4f;
	15'h918: q<=8'h01;
	15'h919: q<=8'hca;
	15'h91a: q<=8'h10;
	15'h91b: q<=8'ha6;
	15'h91c: q<=8'had;
	15'h91d: q<=8'h4f;
	15'h91e: q<=8'h01;
	15'h91f: q<=8'h8d;
	15'h920: q<=8'h50;
	15'h921: q<=8'h01;
	15'h922: q<=8'h60;
	15'h923: q<=8'ha9;
	15'h924: q<=8'hf0;
	15'h925: q<=8'h85;
	15'h926: q<=8'h29;
	15'h927: q<=8'hbd;
	15'h928: q<=8'h03;
	15'h929: q<=8'h02;
	15'h92a: q<=8'h85;
	15'h92b: q<=8'h2a;
	15'h92c: q<=8'h86;
	15'h92d: q<=8'h35;
	15'h92e: q<=8'h20;
	15'h92f: q<=8'ha5;
	15'h930: q<=8'h99;
	15'h931: q<=8'ha6;
	15'h932: q<=8'h35;
	15'h933: q<=8'ha5;
	15'h934: q<=8'h29;
	15'h935: q<=8'hf0;
	15'h936: q<=8'h0e;
	15'h937: q<=8'h20;
	15'h938: q<=8'h4d;
	15'h939: q<=8'h99;
	15'h93a: q<=8'hf0;
	15'h93b: q<=8'h09;
	15'h93c: q<=8'hce;
	15'h93d: q<=8'hab;
	15'h93e: q<=8'h03;
	15'h93f: q<=8'ha9;
	15'h940: q<=8'h00;
	15'h941: q<=8'h9d;
	15'h942: q<=8'h43;
	15'h943: q<=8'h02;
	15'h944: q<=8'h60;
	15'h945: q<=8'ha9;
	15'h946: q<=8'hff;
	15'h947: q<=8'h85;
	15'h948: q<=8'h2f;
	15'h949: q<=8'hfe;
	15'h94a: q<=8'h43;
	15'h94b: q<=8'h02;
	15'h94c: q<=8'h60;
	15'h94d: q<=8'h84;
	15'h94e: q<=8'h36;
	15'h94f: q<=8'hac;
	15'h950: q<=8'h1c;
	15'h951: q<=8'h01;
	15'h952: q<=8'hb9;
	15'h953: q<=8'hdf;
	15'h954: q<=8'h02;
	15'h955: q<=8'hd0;
	15'h956: q<=8'h46;
	15'h957: q<=8'ha5;
	15'h958: q<=8'h29;
	15'h959: q<=8'h99;
	15'h95a: q<=8'hdf;
	15'h95b: q<=8'h02;
	15'h95c: q<=8'ha5;
	15'h95d: q<=8'h2a;
	15'h95e: q<=8'hc9;
	15'h95f: q<=8'h0f;
	15'h960: q<=8'hd0;
	15'h961: q<=8'h0a;
	15'h962: q<=8'h2c;
	15'h963: q<=8'h11;
	15'h964: q<=8'h01;
	15'h965: q<=8'h10;
	15'h966: q<=8'h05;
	15'h967: q<=8'had;
	15'h968: q<=8'hca;
	15'h969: q<=8'h60;
	15'h96a: q<=8'h29;
	15'h96b: q<=8'h0e;
	15'h96c: q<=8'h99;
	15'h96d: q<=8'hb9;
	15'h96e: q<=8'h02;
	15'h96f: q<=8'h18;
	15'h970: q<=8'h69;
	15'h971: q<=8'h01;
	15'h972: q<=8'h29;
	15'h973: q<=8'h0f;
	15'h974: q<=8'h99;
	15'h975: q<=8'hcc;
	15'h976: q<=8'h02;
	15'h977: q<=8'ha9;
	15'h978: q<=8'h00;
	15'h979: q<=8'h99;
	15'h97a: q<=8'ha6;
	15'h97b: q<=8'h02;
	15'h97c: q<=8'ha5;
	15'h97d: q<=8'h2c;
	15'h97e: q<=8'h99;
	15'h97f: q<=8'h8a;
	15'h980: q<=8'h02;
	15'h981: q<=8'ha5;
	15'h982: q<=8'h2d;
	15'h983: q<=8'h99;
	15'h984: q<=8'h91;
	15'h985: q<=8'h02;
	15'h986: q<=8'hee;
	15'h987: q<=8'h08;
	15'h988: q<=8'h01;
	15'h989: q<=8'ha5;
	15'h98a: q<=8'h2b;
	15'h98b: q<=8'h99;
	15'h98c: q<=8'h83;
	15'h98d: q<=8'h02;
	15'h98e: q<=8'ha4;
	15'h98f: q<=8'h36;
	15'h990: q<=8'h29;
	15'h991: q<=8'h07;
	15'h992: q<=8'h86;
	15'h993: q<=8'h36;
	15'h994: q<=8'haa;
	15'h995: q<=8'hfe;
	15'h996: q<=8'h42;
	15'h997: q<=8'h01;
	15'h998: q<=8'ha6;
	15'h999: q<=8'h36;
	15'h99a: q<=8'ha9;
	15'h99b: q<=8'h10;
	15'h99c: q<=8'h60;
	15'h99d: q<=8'h88;
	15'h99e: q<=8'h10;
	15'h99f: q<=8'hb2;
	15'h9a0: q<=8'ha4;
	15'h9a1: q<=8'h36;
	15'h9a2: q<=8'ha9;
	15'h9a3: q<=8'h00;
	15'h9a4: q<=8'h60;
	15'h9a5: q<=8'ha9;
	15'h9a6: q<=8'h00;
	15'h9a7: q<=8'ha2;
	15'h9a8: q<=8'h04;
	15'h9a9: q<=8'h9d;
	15'h9aa: q<=8'h3d;
	15'h9ab: q<=8'h01;
	15'h9ac: q<=8'hca;
	15'h9ad: q<=8'h10;
	15'h9ae: q<=8'hfa;
	15'h9af: q<=8'ha2;
	15'h9b0: q<=8'h04;
	15'h9b1: q<=8'hbd;
	15'h9b2: q<=8'h2e;
	15'h9b3: q<=8'h01;
	15'h9b4: q<=8'h38;
	15'h9b5: q<=8'hfd;
	15'h9b6: q<=8'h42;
	15'h9b7: q<=8'h01;
	15'h9b8: q<=8'h90;
	15'h9b9: q<=8'h03;
	15'h9ba: q<=8'h9d;
	15'h9bb: q<=8'h3d;
	15'h9bc: q<=8'h01;
	15'h9bd: q<=8'hca;
	15'h9be: q<=8'h10;
	15'h9bf: q<=8'hf1;
	15'h9c0: q<=8'hac;
	15'h9c1: q<=8'h1c;
	15'h9c2: q<=8'h01;
	15'h9c3: q<=8'hb9;
	15'h9c4: q<=8'hdf;
	15'h9c5: q<=8'h02;
	15'h9c6: q<=8'hf0;
	15'h9c7: q<=8'h14;
	15'h9c8: q<=8'hb9;
	15'h9c9: q<=8'h8a;
	15'h9ca: q<=8'h02;
	15'h9cb: q<=8'h29;
	15'h9cc: q<=8'h03;
	15'h9cd: q<=8'hf0;
	15'h9ce: q<=8'h0d;
	15'h9cf: q<=8'haa;
	15'h9d0: q<=8'he0;
	15'h9d1: q<=8'h03;
	15'h9d2: q<=8'hd0;
	15'h9d3: q<=8'h02;
	15'h9d4: q<=8'ha2;
	15'h9d5: q<=8'h05;
	15'h9d6: q<=8'hde;
	15'h9d7: q<=8'h3c;
	15'h9d8: q<=8'h01;
	15'h9d9: q<=8'hde;
	15'h9da: q<=8'h3c;
	15'h9db: q<=8'h01;
	15'h9dc: q<=8'h88;
	15'h9dd: q<=8'h10;
	15'h9de: q<=8'he4;
	15'h9df: q<=8'ha2;
	15'h9e0: q<=8'h04;
	15'h9e1: q<=8'had;
	15'h9e2: q<=8'h1c;
	15'h9e3: q<=8'h01;
	15'h9e4: q<=8'h18;
	15'h9e5: q<=8'h69;
	15'h9e6: q<=8'h01;
	15'h9e7: q<=8'h38;
	15'h9e8: q<=8'hfd;
	15'h9e9: q<=8'h42;
	15'h9ea: q<=8'h01;
	15'h9eb: q<=8'hca;
	15'h9ec: q<=8'h10;
	15'h9ed: q<=8'hf9;
	15'h9ee: q<=8'ha2;
	15'h9ef: q<=8'h04;
	15'h9f0: q<=8'hdd;
	15'h9f1: q<=8'h3d;
	15'h9f2: q<=8'h01;
	15'h9f3: q<=8'hb0;
	15'h9f4: q<=8'h03;
	15'h9f5: q<=8'h9d;
	15'h9f6: q<=8'h3d;
	15'h9f7: q<=8'h01;
	15'h9f8: q<=8'hca;
	15'h9f9: q<=8'h10;
	15'h9fa: q<=8'hf5;
	15'h9fb: q<=8'ha2;
	15'h9fc: q<=8'h04;
	15'h9fd: q<=8'ha0;
	15'h9fe: q<=8'h00;
	15'h9ff: q<=8'hbd;
	15'ha00: q<=8'h3d;
	15'ha01: q<=8'h01;
	15'ha02: q<=8'hf0;
	15'ha03: q<=8'h01;
	15'ha04: q<=8'hc8;
	15'ha05: q<=8'hca;
	15'ha06: q<=8'h10;
	15'ha07: q<=8'hf7;
	15'ha08: q<=8'h98;
	15'ha09: q<=8'hf0;
	15'ha0a: q<=8'h77;
	15'ha0b: q<=8'h88;
	15'ha0c: q<=8'hd0;
	15'ha0d: q<=8'h18;
	15'ha0e: q<=8'ha2;
	15'ha0f: q<=8'h04;
	15'ha10: q<=8'hbd;
	15'ha11: q<=8'h3d;
	15'ha12: q<=8'h01;
	15'ha13: q<=8'hf0;
	15'ha14: q<=8'h0b;
	15'ha15: q<=8'hbd;
	15'ha16: q<=8'h29;
	15'ha17: q<=8'h01;
	15'ha18: q<=8'hf0;
	15'ha19: q<=8'h06;
	15'ha1a: q<=8'h20;
	15'ha1b: q<=8'h87;
	15'ha1c: q<=8'h9a;
	15'ha1d: q<=8'hf0;
	15'ha1e: q<=8'h01;
	15'ha1f: q<=8'h60;
	15'ha20: q<=8'hca;
	15'ha21: q<=8'h10;
	15'ha22: q<=8'hed;
	15'ha23: q<=8'hb8;
	15'ha24: q<=8'h50;
	15'ha25: q<=8'h5c;
	15'ha26: q<=8'h84;
	15'ha27: q<=8'h61;
	15'ha28: q<=8'ha2;
	15'ha29: q<=8'h04;
	15'ha2a: q<=8'hbd;
	15'ha2b: q<=8'h3d;
	15'ha2c: q<=8'h01;
	15'ha2d: q<=8'hf0;
	15'ha2e: q<=8'h0e;
	15'ha2f: q<=8'hbd;
	15'ha30: q<=8'h42;
	15'ha31: q<=8'h01;
	15'ha32: q<=8'hdd;
	15'ha33: q<=8'h29;
	15'ha34: q<=8'h01;
	15'ha35: q<=8'hb0;
	15'ha36: q<=8'h06;
	15'ha37: q<=8'h20;
	15'ha38: q<=8'h87;
	15'ha39: q<=8'h9a;
	15'ha3a: q<=8'hf0;
	15'ha3b: q<=8'h01;
	15'ha3c: q<=8'h60;
	15'ha3d: q<=8'hca;
	15'ha3e: q<=8'h10;
	15'ha3f: q<=8'hea;
	15'ha40: q<=8'had;
	15'ha41: q<=8'h40;
	15'ha42: q<=8'h01;
	15'ha43: q<=8'hf0;
	15'ha44: q<=8'h1c;
	15'ha45: q<=8'had;
	15'ha46: q<=8'h3f;
	15'ha47: q<=8'h01;
	15'ha48: q<=8'hf0;
	15'ha49: q<=8'h17;
	15'ha4a: q<=8'ha4;
	15'ha4b: q<=8'h2a;
	15'ha4c: q<=8'hb9;
	15'ha4d: q<=8'hac;
	15'ha4e: q<=8'h03;
	15'ha4f: q<=8'hd0;
	15'ha50: q<=8'h02;
	15'ha51: q<=8'ha9;
	15'ha52: q<=8'hff;
	15'ha53: q<=8'ha2;
	15'ha54: q<=8'h03;
	15'ha55: q<=8'hc9;
	15'ha56: q<=8'hcc;
	15'ha57: q<=8'hb0;
	15'ha58: q<=8'h02;
	15'ha59: q<=8'ha2;
	15'ha5a: q<=8'h02;
	15'ha5b: q<=8'h20;
	15'ha5c: q<=8'h87;
	15'ha5d: q<=8'h9a;
	15'ha5e: q<=8'hf0;
	15'ha5f: q<=8'h01;
	15'ha60: q<=8'h60;
	15'ha61: q<=8'had;
	15'ha62: q<=8'hda;
	15'ha63: q<=8'h60;
	15'ha64: q<=8'h29;
	15'ha65: q<=8'h03;
	15'ha66: q<=8'haa;
	15'ha67: q<=8'he8;
	15'ha68: q<=8'ha0;
	15'ha69: q<=8'h04;
	15'ha6a: q<=8'hbd;
	15'ha6b: q<=8'h29;
	15'ha6c: q<=8'h01;
	15'ha6d: q<=8'hf0;
	15'ha6e: q<=8'h0b;
	15'ha6f: q<=8'hbd;
	15'ha70: q<=8'h3d;
	15'ha71: q<=8'h01;
	15'ha72: q<=8'hf0;
	15'ha73: q<=8'h06;
	15'ha74: q<=8'h20;
	15'ha75: q<=8'h87;
	15'ha76: q<=8'h9a;
	15'ha77: q<=8'hf0;
	15'ha78: q<=8'h01;
	15'ha79: q<=8'h60;
	15'ha7a: q<=8'hca;
	15'ha7b: q<=8'h10;
	15'ha7c: q<=8'h02;
	15'ha7d: q<=8'ha2;
	15'ha7e: q<=8'h04;
	15'ha7f: q<=8'h88;
	15'ha80: q<=8'h10;
	15'ha81: q<=8'he8;
	15'ha82: q<=8'ha9;
	15'ha83: q<=8'h00;
	15'ha84: q<=8'h85;
	15'ha85: q<=8'h29;
	15'ha86: q<=8'h60;
	15'ha87: q<=8'h8a;
	15'ha88: q<=8'h0a;
	15'ha89: q<=8'ha8;
	15'ha8a: q<=8'hb9;
	15'ha8b: q<=8'h94;
	15'ha8c: q<=8'h9a;
	15'ha8d: q<=8'h48;
	15'ha8e: q<=8'hb9;
	15'ha8f: q<=8'h93;
	15'ha90: q<=8'h9a;
	15'ha91: q<=8'h48;
	15'ha92: q<=8'h60;
	15'ha93: q<=8'h9c;
	15'ha94: q<=8'h9a;
	15'ha95: q<=8'ha8;
	15'ha96: q<=8'h9a;
	15'ha97: q<=8'hba;
	15'ha98: q<=8'h9a;
	15'ha99: q<=8'hb6;
	15'ha9a: q<=8'h9a;
	15'ha9b: q<=8'hb2;
	15'ha9c: q<=8'h9a;
	15'ha9d: q<=8'had;
	15'ha9e: q<=8'h02;
	15'ha9f: q<=8'h9b;
	15'haa0: q<=8'h85;
	15'haa1: q<=8'h2c;
	15'haa2: q<=8'had;
	15'haa3: q<=8'h5d;
	15'haa4: q<=8'h01;
	15'haa5: q<=8'ha0;
	15'haa6: q<=8'h00;
	15'haa7: q<=8'hf0;
	15'haa8: q<=8'h4d;
	15'haa9: q<=8'had;
	15'haaa: q<=8'h03;
	15'haab: q<=8'h9b;
	15'haac: q<=8'h0d;
	15'haad: q<=8'h6d;
	15'haae: q<=8'h01;
	15'haaf: q<=8'ha0;
	15'hab0: q<=8'h01;
	15'hab1: q<=8'hd0;
	15'hab2: q<=8'h3e;
	15'hab3: q<=8'ha0;
	15'hab4: q<=8'h04;
	15'hab5: q<=8'hd0;
	15'hab6: q<=8'h37;
	15'hab7: q<=8'ha0;
	15'hab8: q<=8'h03;
	15'hab9: q<=8'hd0;
	15'haba: q<=8'h33;
	15'habb: q<=8'had;
	15'habc: q<=8'hca;
	15'habd: q<=8'h60;
	15'habe: q<=8'h29;
	15'habf: q<=8'h03;
	15'hac0: q<=8'ha8;
	15'hac1: q<=8'ha9;
	15'hac2: q<=8'h04;
	15'hac3: q<=8'h85;
	15'hac4: q<=8'h2b;
	15'hac5: q<=8'h86;
	15'hac6: q<=8'h39;
	15'hac7: q<=8'hc6;
	15'hac8: q<=8'h2b;
	15'hac9: q<=8'h10;
	15'haca: q<=8'h05;
	15'hacb: q<=8'ha6;
	15'hacc: q<=8'h39;
	15'hacd: q<=8'ha9;
	15'hace: q<=8'h00;
	15'hacf: q<=8'h60;
	15'had0: q<=8'h88;
	15'had1: q<=8'h10;
	15'had2: q<=8'h02;
	15'had3: q<=8'ha0;
	15'had4: q<=8'h03;
	15'had5: q<=8'hbe;
	15'had6: q<=8'h49;
	15'had7: q<=8'h01;
	15'had8: q<=8'he0;
	15'had9: q<=8'h03;
	15'hada: q<=8'hd0;
	15'hadb: q<=8'h02;
	15'hadc: q<=8'ha2;
	15'hadd: q<=8'h05;
	15'hade: q<=8'hbd;
	15'hadf: q<=8'h3c;
	15'hae0: q<=8'h01;
	15'hae1: q<=8'hf0;
	15'hae2: q<=8'he4;
	15'hae3: q<=8'ha6;
	15'hae4: q<=8'h39;
	15'hae5: q<=8'hb9;
	15'hae6: q<=8'h49;
	15'hae7: q<=8'h01;
	15'hae8: q<=8'h09;
	15'hae9: q<=8'h40;
	15'haea: q<=8'ha0;
	15'haeb: q<=8'h02;
	15'haec: q<=8'hd0;
	15'haed: q<=8'h03;
	15'haee: q<=8'hb9;
	15'haef: q<=8'h02;
	15'haf0: q<=8'h9b;
	15'haf1: q<=8'h85;
	15'haf2: q<=8'h2c;
	15'haf3: q<=8'hb9;
	15'haf4: q<=8'hfd;
	15'haf5: q<=8'h9a;
	15'haf6: q<=8'h84;
	15'haf7: q<=8'h2b;
	15'haf8: q<=8'h85;
	15'haf9: q<=8'h2d;
	15'hafa: q<=8'ha5;
	15'hafb: q<=8'h29;
	15'hafc: q<=8'h60;
	15'hafd: q<=8'h07;
	15'hafe: q<=8'h72;
	15'haff: q<=8'h07;
	15'hb00: q<=8'h00;
	15'hb01: q<=8'h61;
	15'hb02: q<=8'h40;
	15'hb03: q<=8'h00;
	15'hb04: q<=8'h41;
	15'hb05: q<=8'h40;
	15'hb06: q<=8'h00;
	15'hb07: q<=8'h84;
	15'hb08: q<=8'h36;
	15'hb09: q<=8'ha5;
	15'hb0a: q<=8'h29;
	15'hb0b: q<=8'hc9;
	15'hb0c: q<=8'h20;
	15'hb0d: q<=8'ha5;
	15'hb0e: q<=8'h2b;
	15'hb0f: q<=8'hb0;
	15'hb10: q<=8'h07;
	15'hb11: q<=8'ha8;
	15'hb12: q<=8'h20;
	15'hb13: q<=8'hee;
	15'hb14: q<=8'h9a;
	15'hb15: q<=8'hb8;
	15'hb16: q<=8'h50;
	15'hb17: q<=8'h03;
	15'hb18: q<=8'h20;
	15'hb19: q<=8'h88;
	15'hb1a: q<=8'h9a;
	15'hb1b: q<=8'ha4;
	15'hb1c: q<=8'h36;
	15'hb1d: q<=8'h60;
	15'hb1e: q<=8'had;
	15'hb1f: q<=8'h01;
	15'hb20: q<=8'h02;
	15'hb21: q<=8'h30;
	15'hb22: q<=8'h33;
	15'hb23: q<=8'hae;
	15'hb24: q<=8'h1c;
	15'hb25: q<=8'h01;
	15'hb26: q<=8'h86;
	15'hb27: q<=8'h37;
	15'hb28: q<=8'ha6;
	15'hb29: q<=8'h37;
	15'hb2a: q<=8'hbd;
	15'hb2b: q<=8'hdf;
	15'hb2c: q<=8'h02;
	15'hb2d: q<=8'hf0;
	15'hb2e: q<=8'h23;
	15'hb2f: q<=8'ha9;
	15'hb30: q<=8'h01;
	15'hb31: q<=8'h8d;
	15'hb32: q<=8'h0a;
	15'hb33: q<=8'h01;
	15'hb34: q<=8'hbd;
	15'hb35: q<=8'h91;
	15'hb36: q<=8'h02;
	15'hb37: q<=8'h8d;
	15'hb38: q<=8'h0b;
	15'hb39: q<=8'h01;
	15'hb3a: q<=8'had;
	15'hb3b: q<=8'h0b;
	15'hb3c: q<=8'h01;
	15'hb3d: q<=8'ha8;
	15'hb3e: q<=8'hb9;
	15'hb3f: q<=8'hf7;
	15'hb40: q<=8'ha0;
	15'hb41: q<=8'h20;
	15'hb42: q<=8'h98;
	15'hb43: q<=8'h9b;
	15'hb44: q<=8'hee;
	15'hb45: q<=8'h0b;
	15'hb46: q<=8'h01;
	15'hb47: q<=8'had;
	15'hb48: q<=8'h0a;
	15'hb49: q<=8'h01;
	15'hb4a: q<=8'hd0;
	15'hb4b: q<=8'hee;
	15'hb4c: q<=8'had;
	15'hb4d: q<=8'h0b;
	15'hb4e: q<=8'h01;
	15'hb4f: q<=8'h9d;
	15'hb50: q<=8'h91;
	15'hb51: q<=8'h02;
	15'hb52: q<=8'hc6;
	15'hb53: q<=8'h37;
	15'hb54: q<=8'h10;
	15'hb55: q<=8'hd2;
	15'hb56: q<=8'had;
	15'hb57: q<=8'h48;
	15'hb58: q<=8'h01;
	15'hb59: q<=8'h18;
	15'hb5a: q<=8'h6d;
	15'hb5b: q<=8'h47;
	15'hb5c: q<=8'h01;
	15'hb5d: q<=8'ha8;
	15'hb5e: q<=8'h4d;
	15'hb5f: q<=8'h48;
	15'hb60: q<=8'h01;
	15'hb61: q<=8'h8c;
	15'hb62: q<=8'h48;
	15'hb63: q<=8'h01;
	15'hb64: q<=8'h10;
	15'hb65: q<=8'h16;
	15'hb66: q<=8'h98;
	15'hb67: q<=8'h10;
	15'hb68: q<=8'h06;
	15'hb69: q<=8'h20;
	15'hb6a: q<=8'h06;
	15'hb6b: q<=8'hcd;
	15'hb6c: q<=8'hb8;
	15'hb6d: q<=8'h50;
	15'hb6e: q<=8'h0d;
	15'hb6f: q<=8'had;
	15'hb70: q<=8'h43;
	15'hb71: q<=8'h01;
	15'hb72: q<=8'hf0;
	15'hb73: q<=8'h08;
	15'hb74: q<=8'had;
	15'hb75: q<=8'h01;
	15'hb76: q<=8'h02;
	15'hb77: q<=8'h30;
	15'hb78: q<=8'h03;
	15'hb79: q<=8'h20;
	15'hb7a: q<=8'h02;
	15'hb7b: q<=8'hcd;
	15'hb7c: q<=8'had;
	15'hb7d: q<=8'h48;
	15'hb7e: q<=8'h01;
	15'hb7f: q<=8'h30;
	15'hb80: q<=8'h07;
	15'hb81: q<=8'hc9;
	15'hb82: q<=8'h0f;
	15'hb83: q<=8'hb0;
	15'hb84: q<=8'h07;
	15'hb85: q<=8'hb8;
	15'hb86: q<=8'h50;
	15'hb87: q<=8'h0f;
	15'hb88: q<=8'hc9;
	15'hb89: q<=8'hc1;
	15'hb8a: q<=8'hb0;
	15'hb8b: q<=8'h0b;
	15'hb8c: q<=8'had;
	15'hb8d: q<=8'h47;
	15'hb8e: q<=8'h01;
	15'hb8f: q<=8'h49;
	15'hb90: q<=8'hff;
	15'hb91: q<=8'h18;
	15'hb92: q<=8'h69;
	15'hb93: q<=8'h01;
	15'hb94: q<=8'h8d;
	15'hb95: q<=8'h47;
	15'hb96: q<=8'h01;
	15'hb97: q<=8'h60;
	15'hb98: q<=8'ha8;
	15'hb99: q<=8'hb9;
	15'hb9a: q<=8'ha3;
	15'hb9b: q<=8'h9b;
	15'hb9c: q<=8'h48;
	15'hb9d: q<=8'hb9;
	15'hb9e: q<=8'ha2;
	15'hb9f: q<=8'h9b;
	15'hba0: q<=8'h48;
	15'hba1: q<=8'h60;
	15'hba2: q<=8'hc9;
	15'hba3: q<=8'h9b;
	15'hba4: q<=8'hcf;
	15'hba5: q<=8'h9b;
	15'hba6: q<=8'hed;
	15'hba7: q<=8'h9b;
	15'hba8: q<=8'h16;
	15'hba9: q<=8'h9c;
	15'hbaa: q<=8'h0b;
	15'hbab: q<=8'h9c;
	15'hbac: q<=8'hce;
	15'hbad: q<=8'h9b;
	15'hbae: q<=8'h57;
	15'hbaf: q<=8'h9c;
	15'hbb0: q<=8'hc3;
	15'hbb1: q<=8'h9f;
	15'hbb2: q<=8'hdc;
	15'hbb3: q<=8'h9b;
	15'hbb4: q<=8'h5b;
	15'hbb5: q<=8'h9e;
	15'hbb6: q<=8'h81;
	15'hbb7: q<=8'h9d;
	15'hbb8: q<=8'h4e;
	15'hbb9: q<=8'h9c;
	15'hbba: q<=8'h2e;
	15'hbbb: q<=8'h9e;
	15'hbbc: q<=8'hf9;
	15'hbbd: q<=8'h9b;
	15'hbbe: q<=8'h20;
	15'hbbf: q<=8'h9c;
	15'hbc0: q<=8'hf0;
	15'hbc1: q<=8'h9e;
	15'hbc2: q<=8'h47;
	15'hbc3: q<=8'h9e;
	15'hbc4: q<=8'hb5;
	15'hbc5: q<=8'h9c;
	15'hbc6: q<=8'h66;
	15'hbc7: q<=8'h9d;
	15'hbc8: q<=8'h3a;
	15'hbc9: q<=8'h9c;
	15'hbca: q<=8'ha9;
	15'hbcb: q<=8'h00;
	15'hbcc: q<=8'h8d;
	15'hbcd: q<=8'h0a;
	15'hbce: q<=8'h01;
	15'hbcf: q<=8'h60;
	15'hbd0: q<=8'hee;
	15'hbd1: q<=8'h0b;
	15'hbd2: q<=8'h01;
	15'hbd3: q<=8'hac;
	15'hbd4: q<=8'h0b;
	15'hbd5: q<=8'h01;
	15'hbd6: q<=8'hb9;
	15'hbd7: q<=8'hf7;
	15'hbd8: q<=8'ha0;
	15'hbd9: q<=8'h9d;
	15'hbda: q<=8'h98;
	15'hbdb: q<=8'h02;
	15'hbdc: q<=8'h60;
	15'hbdd: q<=8'hee;
	15'hbde: q<=8'h0b;
	15'hbdf: q<=8'h01;
	15'hbe0: q<=8'hac;
	15'hbe1: q<=8'h0b;
	15'hbe2: q<=8'h01;
	15'hbe3: q<=8'hb9;
	15'hbe4: q<=8'hf7;
	15'hbe5: q<=8'ha0;
	15'hbe6: q<=8'ha8;
	15'hbe7: q<=8'hb9;
	15'hbe8: q<=8'h00;
	15'hbe9: q<=8'h00;
	15'hbea: q<=8'h9d;
	15'hbeb: q<=8'h98;
	15'hbec: q<=8'h02;
	15'hbed: q<=8'h60;
	15'hbee: q<=8'had;
	15'hbef: q<=8'h0c;
	15'hbf0: q<=8'h01;
	15'hbf1: q<=8'hd0;
	15'hbf2: q<=8'h06;
	15'hbf3: q<=8'hee;
	15'hbf4: q<=8'h0b;
	15'hbf5: q<=8'h01;
	15'hbf6: q<=8'hee;
	15'hbf7: q<=8'h0b;
	15'hbf8: q<=8'h01;
	15'hbf9: q<=8'h60;
	15'hbfa: q<=8'hee;
	15'hbfb: q<=8'h0b;
	15'hbfc: q<=8'h01;
	15'hbfd: q<=8'had;
	15'hbfe: q<=8'h0c;
	15'hbff: q<=8'h01;
	15'hc00: q<=8'hd0;
	15'hc01: q<=8'h09;
	15'hc02: q<=8'hac;
	15'hc03: q<=8'h0b;
	15'hc04: q<=8'h01;
	15'hc05: q<=8'hb9;
	15'hc06: q<=8'hf7;
	15'hc07: q<=8'ha0;
	15'hc08: q<=8'h8d;
	15'hc09: q<=8'h0b;
	15'hc0a: q<=8'h01;
	15'hc0b: q<=8'h60;
	15'hc0c: q<=8'hde;
	15'hc0d: q<=8'h98;
	15'hc0e: q<=8'h02;
	15'hc0f: q<=8'hd0;
	15'hc10: q<=8'h06;
	15'hc11: q<=8'hee;
	15'hc12: q<=8'h0b;
	15'hc13: q<=8'h01;
	15'hc14: q<=8'hb8;
	15'hc15: q<=8'h50;
	15'hc16: q<=8'h09;
	15'hc17: q<=8'hac;
	15'hc18: q<=8'h0b;
	15'hc19: q<=8'h01;
	15'hc1a: q<=8'hb9;
	15'hc1b: q<=8'hf8;
	15'hc1c: q<=8'ha0;
	15'hc1d: q<=8'h8d;
	15'hc1e: q<=8'h0b;
	15'hc1f: q<=8'h01;
	15'hc20: q<=8'h60;
	15'hc21: q<=8'hbc;
	15'hc22: q<=8'hb9;
	15'hc23: q<=8'h02;
	15'hc24: q<=8'hb9;
	15'hc25: q<=8'hac;
	15'hc26: q<=8'h03;
	15'hc27: q<=8'hd0;
	15'hc28: q<=8'h02;
	15'hc29: q<=8'ha9;
	15'hc2a: q<=8'hff;
	15'hc2b: q<=8'hdd;
	15'hc2c: q<=8'hdf;
	15'hc2d: q<=8'h02;
	15'hc2e: q<=8'hb0;
	15'hc2f: q<=8'h05;
	15'hc30: q<=8'ha9;
	15'hc31: q<=8'h00;
	15'hc32: q<=8'hb8;
	15'hc33: q<=8'h50;
	15'hc34: q<=8'h02;
	15'hc35: q<=8'ha9;
	15'hc36: q<=8'h01;
	15'hc37: q<=8'h8d;
	15'hc38: q<=8'h0c;
	15'hc39: q<=8'h01;
	15'hc3a: q<=8'h60;
	15'hc3b: q<=8'had;
	15'hc3c: q<=8'h47;
	15'hc3d: q<=8'h01;
	15'hc3e: q<=8'h0a;
	15'hc3f: q<=8'h0a;
	15'hc40: q<=8'h18;
	15'hc41: q<=8'h6d;
	15'hc42: q<=8'h48;
	15'hc43: q<=8'h01;
	15'hc44: q<=8'h2d;
	15'hc45: q<=8'h48;
	15'hc46: q<=8'h01;
	15'hc47: q<=8'h29;
	15'hc48: q<=8'h80;
	15'hc49: q<=8'h49;
	15'hc4a: q<=8'h80;
	15'hc4b: q<=8'h8d;
	15'hc4c: q<=8'h0c;
	15'hc4d: q<=8'h01;
	15'hc4e: q<=8'h60;
	15'hc4f: q<=8'hbd;
	15'hc50: q<=8'h83;
	15'hc51: q<=8'h02;
	15'hc52: q<=8'h49;
	15'hc53: q<=8'h40;
	15'hc54: q<=8'h9d;
	15'hc55: q<=8'h83;
	15'hc56: q<=8'h02;
	15'hc57: q<=8'h60;
	15'hc58: q<=8'hbd;
	15'hc59: q<=8'h83;
	15'hc5a: q<=8'h02;
	15'hc5b: q<=8'h29;
	15'hc5c: q<=8'h07;
	15'hc5d: q<=8'ha8;
	15'hc5e: q<=8'hbd;
	15'hc5f: q<=8'h8a;
	15'hc60: q<=8'h02;
	15'hc61: q<=8'h30;
	15'hc62: q<=8'h36;
	15'hc63: q<=8'hbd;
	15'hc64: q<=8'h9f;
	15'hc65: q<=8'h02;
	15'hc66: q<=8'h18;
	15'hc67: q<=8'h79;
	15'hc68: q<=8'h60;
	15'hc69: q<=8'h01;
	15'hc6a: q<=8'h9d;
	15'hc6b: q<=8'h9f;
	15'hc6c: q<=8'h02;
	15'hc6d: q<=8'hbd;
	15'hc6e: q<=8'hdf;
	15'hc6f: q<=8'h02;
	15'hc70: q<=8'h79;
	15'hc71: q<=8'h65;
	15'hc72: q<=8'h01;
	15'hc73: q<=8'h9d;
	15'hc74: q<=8'hdf;
	15'hc75: q<=8'h02;
	15'hc76: q<=8'hcd;
	15'hc77: q<=8'h02;
	15'hc78: q<=8'h02;
	15'hc79: q<=8'hf0;
	15'hc7a: q<=8'h02;
	15'hc7b: q<=8'hb0;
	15'hc7c: q<=8'h06;
	15'hc7d: q<=8'h20;
	15'hc7e: q<=8'h06;
	15'hc7f: q<=8'h9d;
	15'hc80: q<=8'hb8;
	15'hc81: q<=8'h50;
	15'hc82: q<=8'h13;
	15'hc83: q<=8'hc9;
	15'hc84: q<=8'h20;
	15'hc85: q<=8'hb0;
	15'hc86: q<=8'h0f;
	15'hc87: q<=8'hbd;
	15'hc88: q<=8'h8a;
	15'hc89: q<=8'h02;
	15'hc8a: q<=8'h29;
	15'hc8b: q<=8'h03;
	15'hc8c: q<=8'hf0;
	15'hc8d: q<=8'h08;
	15'hc8e: q<=8'h8a;
	15'hc8f: q<=8'h48;
	15'hc90: q<=8'ha8;
	15'hc91: q<=8'h20;
	15'hc92: q<=8'h6f;
	15'hc93: q<=8'ha0;
	15'hc94: q<=8'h68;
	15'hc95: q<=8'haa;
	15'hc96: q<=8'hb8;
	15'hc97: q<=8'h50;
	15'hc98: q<=8'h1c;
	15'hc99: q<=8'hbd;
	15'hc9a: q<=8'h9f;
	15'hc9b: q<=8'h02;
	15'hc9c: q<=8'h38;
	15'hc9d: q<=8'hf9;
	15'hc9e: q<=8'h60;
	15'hc9f: q<=8'h01;
	15'hca0: q<=8'h9d;
	15'hca1: q<=8'h9f;
	15'hca2: q<=8'h02;
	15'hca3: q<=8'hbd;
	15'hca4: q<=8'hdf;
	15'hca5: q<=8'h02;
	15'hca6: q<=8'hf9;
	15'hca7: q<=8'h65;
	15'hca8: q<=8'h01;
	15'hca9: q<=8'h9d;
	15'hcaa: q<=8'hdf;
	15'hcab: q<=8'h02;
	15'hcac: q<=8'hc9;
	15'hcad: q<=8'hf0;
	15'hcae: q<=8'h90;
	15'hcaf: q<=8'h05;
	15'hcb0: q<=8'ha9;
	15'hcb1: q<=8'hf2;
	15'hcb2: q<=8'h9d;
	15'hcb3: q<=8'hdf;
	15'hcb4: q<=8'h02;
	15'hcb5: q<=8'h60;
	15'hcb6: q<=8'ha0;
	15'hcb7: q<=8'h01;
	15'hcb8: q<=8'hbd;
	15'hcb9: q<=8'h8a;
	15'hcba: q<=8'h02;
	15'hcbb: q<=8'h30;
	15'hcbc: q<=8'h10;
	15'hcbd: q<=8'hbd;
	15'hcbe: q<=8'hdf;
	15'hcbf: q<=8'h02;
	15'hcc0: q<=8'hcd;
	15'hcc1: q<=8'h57;
	15'hcc2: q<=8'h01;
	15'hcc3: q<=8'h90;
	15'hcc4: q<=8'h02;
	15'hcc5: q<=8'ha0;
	15'hcc6: q<=8'h00;
	15'hcc7: q<=8'h20;
	15'hcc8: q<=8'h63;
	15'hcc9: q<=8'h9c;
	15'hcca: q<=8'hb8;
	15'hccb: q<=8'h50;
	15'hccc: q<=8'h17;
	15'hccd: q<=8'h20;
	15'hcce: q<=8'h99;
	15'hccf: q<=8'h9c;
	15'hcd0: q<=8'hac;
	15'hcd1: q<=8'hab;
	15'hcd2: q<=8'h03;
	15'hcd3: q<=8'hd0;
	15'hcd4: q<=8'h02;
	15'hcd5: q<=8'ha9;
	15'hcd6: q<=8'hff;
	15'hcd7: q<=8'hcd;
	15'hcd8: q<=8'h57;
	15'hcd9: q<=8'h01;
	15'hcda: q<=8'h90;
	15'hcdb: q<=8'h08;
	15'hcdc: q<=8'hbd;
	15'hcdd: q<=8'h8a;
	15'hcde: q<=8'h02;
	15'hcdf: q<=8'h49;
	15'hce0: q<=8'h80;
	15'hce1: q<=8'h9d;
	15'hce2: q<=8'h8a;
	15'hce3: q<=8'h02;
	15'hce4: q<=8'had;
	15'hce5: q<=8'h48;
	15'hce6: q<=8'h01;
	15'hce7: q<=8'h30;
	15'hce8: q<=8'h1b;
	15'hce9: q<=8'hbd;
	15'hcea: q<=8'hdf;
	15'hceb: q<=8'h02;
	15'hcec: q<=8'hcd;
	15'hced: q<=8'h57;
	15'hcee: q<=8'h01;
	15'hcef: q<=8'hb0;
	15'hcf0: q<=8'h13;
	15'hcf1: q<=8'had;
	15'hcf2: q<=8'h00;
	15'hcf3: q<=8'h02;
	15'hcf4: q<=8'hdd;
	15'hcf5: q<=8'hb9;
	15'hcf6: q<=8'h02;
	15'hcf7: q<=8'hd0;
	15'hcf8: q<=8'h0b;
	15'hcf9: q<=8'had;
	15'hcfa: q<=8'h01;
	15'hcfb: q<=8'h02;
	15'hcfc: q<=8'hdd;
	15'hcfd: q<=8'hcc;
	15'hcfe: q<=8'h02;
	15'hcff: q<=8'hd0;
	15'hd00: q<=8'h03;
	15'hd01: q<=8'h20;
	15'hd02: q<=8'h47;
	15'hd03: q<=8'ha3;
	15'hd04: q<=8'h60;
	15'hd05: q<=8'h16;
	15'hd06: q<=8'had;
	15'hd07: q<=8'h02;
	15'hd08: q<=8'h02;
	15'hd09: q<=8'h9d;
	15'hd0a: q<=8'hdf;
	15'hd0b: q<=8'h02;
	15'hd0c: q<=8'hbd;
	15'hd0d: q<=8'h83;
	15'hd0e: q<=8'h02;
	15'hd0f: q<=8'h29;
	15'hd10: q<=8'h07;
	15'hd11: q<=8'hc9;
	15'hd12: q<=8'h01;
	15'hd13: q<=8'hd0;
	15'hd14: q<=8'h0e;
	15'hd15: q<=8'had;
	15'hd16: q<=8'hab;
	15'hd17: q<=8'h03;
	15'hd18: q<=8'hf0;
	15'hd19: q<=8'h09;
	15'hd1a: q<=8'hbd;
	15'hd1b: q<=8'h8a;
	15'hd1c: q<=8'h02;
	15'hd1d: q<=8'h49;
	15'hd1e: q<=8'h80;
	15'hd1f: q<=8'h9d;
	15'hd20: q<=8'h8a;
	15'hd21: q<=8'h02;
	15'hd22: q<=8'h60;
	15'hd23: q<=8'hbd;
	15'hd24: q<=8'h83;
	15'hd25: q<=8'h02;
	15'hd26: q<=8'h10;
	15'hd27: q<=8'h04;
	15'hd28: q<=8'hfe;
	15'hd29: q<=8'hdf;
	15'hd2a: q<=8'h02;
	15'hd2b: q<=8'h60;
	15'hd2c: q<=8'hce;
	15'hd2d: q<=8'h08;
	15'hd2e: q<=8'h01;
	15'hd2f: q<=8'had;
	15'hd30: q<=8'h09;
	15'hd31: q<=8'h01;
	15'hd32: q<=8'hc9;
	15'hd33: q<=8'h01;
	15'hd34: q<=8'hf0;
	15'hd35: q<=8'h06;
	15'hd36: q<=8'h20;
	15'hd37: q<=8'h67;
	15'hd38: q<=8'h9d;
	15'hd39: q<=8'hb8;
	15'hd3a: q<=8'h50;
	15'hd3b: q<=8'h22;
	15'hd3c: q<=8'ha0;
	15'hd3d: q<=8'h06;
	15'hd3e: q<=8'hb9;
	15'hd3f: q<=8'hdf;
	15'hd40: q<=8'h02;
	15'hd41: q<=8'hf0;
	15'hd42: q<=8'h0e;
	15'hd43: q<=8'h84;
	15'hd44: q<=8'h38;
	15'hd45: q<=8'he4;
	15'hd46: q<=8'h38;
	15'hd47: q<=8'hf0;
	15'hd48: q<=8'h08;
	15'hd49: q<=8'hb9;
	15'hd4a: q<=8'hdf;
	15'hd4b: q<=8'h02;
	15'hd4c: q<=8'hcd;
	15'hd4d: q<=8'h02;
	15'hd4e: q<=8'h02;
	15'hd4f: q<=8'hf0;
	15'hd50: q<=8'h03;
	15'hd51: q<=8'h88;
	15'hd52: q<=8'h10;
	15'hd53: q<=8'hea;
	15'hd54: q<=8'hb9;
	15'hd55: q<=8'h83;
	15'hd56: q<=8'h02;
	15'hd57: q<=8'h29;
	15'hd58: q<=8'h40;
	15'hd59: q<=8'h49;
	15'hd5a: q<=8'h40;
	15'hd5b: q<=8'h9d;
	15'hd5c: q<=8'h83;
	15'hd5d: q<=8'h02;
	15'hd5e: q<=8'ha9;
	15'hd5f: q<=8'h41;
	15'hd60: q<=8'h8d;
	15'hd61: q<=8'h0b;
	15'hd62: q<=8'h01;
	15'hd63: q<=8'hee;
	15'hd64: q<=8'h09;
	15'hd65: q<=8'h01;
	15'hd66: q<=8'h60;
	15'hd67: q<=8'hbd;
	15'hd68: q<=8'hb9;
	15'hd69: q<=8'h02;
	15'hd6a: q<=8'ha8;
	15'hd6b: q<=8'had;
	15'hd6c: q<=8'h00;
	15'hd6d: q<=8'h02;
	15'hd6e: q<=8'h20;
	15'hd6f: q<=8'ha6;
	15'hd70: q<=8'ha7;
	15'hd71: q<=8'h0a;
	15'hd72: q<=8'hbd;
	15'hd73: q<=8'h83;
	15'hd74: q<=8'h02;
	15'hd75: q<=8'hb0;
	15'hd76: q<=8'h05;
	15'hd77: q<=8'h09;
	15'hd78: q<=8'h40;
	15'hd79: q<=8'hb8;
	15'hd7a: q<=8'h50;
	15'hd7b: q<=8'h02;
	15'hd7c: q<=8'h29;
	15'hd7d: q<=8'hbf;
	15'hd7e: q<=8'h9d;
	15'hd7f: q<=8'h83;
	15'hd80: q<=8'h02;
	15'hd81: q<=8'h60;
	15'hd82: q<=8'hbc;
	15'hd83: q<=8'hcc;
	15'hd84: q<=8'h02;
	15'hd85: q<=8'hbd;
	15'hd86: q<=8'h83;
	15'hd87: q<=8'h02;
	15'hd88: q<=8'h29;
	15'hd89: q<=8'h40;
	15'hd8a: q<=8'hd0;
	15'hd8b: q<=8'h04;
	15'hd8c: q<=8'hc8;
	15'hd8d: q<=8'hb8;
	15'hd8e: q<=8'h50;
	15'hd8f: q<=8'h01;
	15'hd90: q<=8'h88;
	15'hd91: q<=8'h98;
	15'hd92: q<=8'h29;
	15'hd93: q<=8'h0f;
	15'hd94: q<=8'h09;
	15'hd95: q<=8'h80;
	15'hd96: q<=8'h9d;
	15'hd97: q<=8'hcc;
	15'hd98: q<=8'h02;
	15'hd99: q<=8'hbd;
	15'hd9a: q<=8'h83;
	15'hd9b: q<=8'h02;
	15'hd9c: q<=8'h29;
	15'hd9d: q<=8'h07;
	15'hd9e: q<=8'hc9;
	15'hd9f: q<=8'h04;
	15'hda0: q<=8'hd0;
	15'hda1: q<=8'h4c;
	15'hda2: q<=8'hbd;
	15'hda3: q<=8'hcc;
	15'hda4: q<=8'h02;
	15'hda5: q<=8'h29;
	15'hda6: q<=8'h07;
	15'hda7: q<=8'hd0;
	15'hda8: q<=8'h42;
	15'hda9: q<=8'hbd;
	15'hdaa: q<=8'hcc;
	15'hdab: q<=8'h02;
	15'hdac: q<=8'h29;
	15'hdad: q<=8'h08;
	15'hdae: q<=8'hf0;
	15'hdaf: q<=8'h0b;
	15'hdb0: q<=8'hbd;
	15'hdb1: q<=8'hb9;
	15'hdb2: q<=8'h02;
	15'hdb3: q<=8'h18;
	15'hdb4: q<=8'h69;
	15'hdb5: q<=8'h01;
	15'hdb6: q<=8'h29;
	15'hdb7: q<=8'h0f;
	15'hdb8: q<=8'h9d;
	15'hdb9: q<=8'hb9;
	15'hdba: q<=8'h02;
	15'hdbb: q<=8'hbd;
	15'hdbc: q<=8'h83;
	15'hdbd: q<=8'h02;
	15'hdbe: q<=8'h29;
	15'hdbf: q<=8'h7f;
	15'hdc0: q<=8'h9d;
	15'hdc1: q<=8'h83;
	15'hdc2: q<=8'h02;
	15'hdc3: q<=8'ha9;
	15'hdc4: q<=8'h20;
	15'hdc5: q<=8'h9d;
	15'hdc6: q<=8'hcc;
	15'hdc7: q<=8'h02;
	15'hdc8: q<=8'hbd;
	15'hdc9: q<=8'h8a;
	15'hdca: q<=8'h02;
	15'hdcb: q<=8'h49;
	15'hdcc: q<=8'h80;
	15'hdcd: q<=8'h9d;
	15'hdce: q<=8'h8a;
	15'hdcf: q<=8'h02;
	15'hdd0: q<=8'had;
	15'hdd1: q<=8'hab;
	15'hdd2: q<=8'h03;
	15'hdd3: q<=8'hd0;
	15'hdd4: q<=8'h16;
	15'hdd5: q<=8'hbd;
	15'hdd6: q<=8'hdf;
	15'hdd7: q<=8'h02;
	15'hdd8: q<=8'hcd;
	15'hdd9: q<=8'h02;
	15'hdda: q<=8'h02;
	15'hddb: q<=8'hd0;
	15'hddc: q<=8'h06;
	15'hddd: q<=8'h20;
	15'hdde: q<=8'h81;
	15'hddf: q<=8'h9f;
	15'hde0: q<=8'hb8;
	15'hde1: q<=8'h50;
	15'hde2: q<=8'h08;
	15'hde3: q<=8'hbd;
	15'hde4: q<=8'h8a;
	15'hde5: q<=8'h02;
	15'hde6: q<=8'h29;
	15'hde7: q<=8'h80;
	15'hde8: q<=8'h9d;
	15'hde9: q<=8'h8a;
	15'hdea: q<=8'h02;
	15'hdeb: q<=8'hb8;
	15'hdec: q<=8'h50;
	15'hded: q<=8'h38;
	15'hdee: q<=8'hbc;
	15'hdef: q<=8'hb9;
	15'hdf0: q<=8'h02;
	15'hdf1: q<=8'hbd;
	15'hdf2: q<=8'h83;
	15'hdf3: q<=8'h02;
	15'hdf4: q<=8'h49;
	15'hdf5: q<=8'h40;
	15'hdf6: q<=8'h20;
	15'hdf7: q<=8'hd7;
	15'hdf8: q<=8'h9e;
	15'hdf9: q<=8'hdd;
	15'hdfa: q<=8'hcc;
	15'hdfb: q<=8'h02;
	15'hdfc: q<=8'hd0;
	15'hdfd: q<=8'h28;
	15'hdfe: q<=8'hbd;
	15'hdff: q<=8'h83;
	15'he00: q<=8'h02;
	15'he01: q<=8'h29;
	15'he02: q<=8'h7f;
	15'he03: q<=8'h9d;
	15'he04: q<=8'h83;
	15'he05: q<=8'h02;
	15'he06: q<=8'h29;
	15'he07: q<=8'h40;
	15'he08: q<=8'hd0;
	15'he09: q<=8'h11;
	15'he0a: q<=8'hbd;
	15'he0b: q<=8'hb9;
	15'he0c: q<=8'h02;
	15'he0d: q<=8'h9d;
	15'he0e: q<=8'hcc;
	15'he0f: q<=8'h02;
	15'he10: q<=8'h38;
	15'he11: q<=8'he9;
	15'he12: q<=8'h01;
	15'he13: q<=8'h29;
	15'he14: q<=8'h0f;
	15'he15: q<=8'h9d;
	15'he16: q<=8'hb9;
	15'he17: q<=8'h02;
	15'he18: q<=8'hb8;
	15'he19: q<=8'h50;
	15'he1a: q<=8'h0b;
	15'he1b: q<=8'hbd;
	15'he1c: q<=8'hb9;
	15'he1d: q<=8'h02;
	15'he1e: q<=8'h18;
	15'he1f: q<=8'h69;
	15'he20: q<=8'h01;
	15'he21: q<=8'h29;
	15'he22: q<=8'h0f;
	15'he23: q<=8'h9d;
	15'he24: q<=8'hcc;
	15'he25: q<=8'h02;
	15'he26: q<=8'hbd;
	15'he27: q<=8'h83;
	15'he28: q<=8'h02;
	15'he29: q<=8'h29;
	15'he2a: q<=8'h80;
	15'he2b: q<=8'h8d;
	15'he2c: q<=8'h0c;
	15'he2d: q<=8'h01;
	15'he2e: q<=8'h60;
	15'he2f: q<=8'hbd;
	15'he30: q<=8'h83;
	15'he31: q<=8'h02;
	15'he32: q<=8'h30;
	15'he33: q<=8'h13;
	15'he34: q<=8'hbd;
	15'he35: q<=8'hb9;
	15'he36: q<=8'h02;
	15'he37: q<=8'hcd;
	15'he38: q<=8'h00;
	15'he39: q<=8'h02;
	15'he3a: q<=8'hd0;
	15'he3b: q<=8'h0b;
	15'he3c: q<=8'hbd;
	15'he3d: q<=8'hcc;
	15'he3e: q<=8'h02;
	15'he3f: q<=8'hcd;
	15'he40: q<=8'h01;
	15'he41: q<=8'h02;
	15'he42: q<=8'hd0;
	15'he43: q<=8'h03;
	15'he44: q<=8'h20;
	15'he45: q<=8'h3a;
	15'he46: q<=8'ha3;
	15'he47: q<=8'h60;
	15'he48: q<=8'hbd;
	15'he49: q<=8'hdf;
	15'he4a: q<=8'h02;
	15'he4b: q<=8'hcd;
	15'he4c: q<=8'h02;
	15'he4d: q<=8'h02;
	15'he4e: q<=8'hd0;
	15'he4f: q<=8'h0b;
	15'he50: q<=8'hbd;
	15'he51: q<=8'hb9;
	15'he52: q<=8'h02;
	15'he53: q<=8'hcd;
	15'he54: q<=8'h00;
	15'he55: q<=8'h02;
	15'he56: q<=8'hd0;
	15'he57: q<=8'h03;
	15'he58: q<=8'h20;
	15'he59: q<=8'h43;
	15'he5a: q<=8'ha3;
	15'he5b: q<=8'h60;
	15'he5c: q<=8'h20;
	15'he5d: q<=8'hab;
	15'he5e: q<=8'h9e;
	15'he5f: q<=8'hbd;
	15'he60: q<=8'h83;
	15'he61: q<=8'h02;
	15'he62: q<=8'h09;
	15'he63: q<=8'h80;
	15'he64: q<=8'h9d;
	15'he65: q<=8'h83;
	15'he66: q<=8'h02;
	15'he67: q<=8'h29;
	15'he68: q<=8'h07;
	15'he69: q<=8'hc9;
	15'he6a: q<=8'h04;
	15'he6b: q<=8'hd0;
	15'he6c: q<=8'h1f;
	15'he6d: q<=8'hbd;
	15'he6e: q<=8'h83;
	15'he6f: q<=8'h02;
	15'he70: q<=8'h29;
	15'he71: q<=8'h40;
	15'he72: q<=8'hd0;
	15'he73: q<=8'h05;
	15'he74: q<=8'ha9;
	15'he75: q<=8'h81;
	15'he76: q<=8'hb8;
	15'he77: q<=8'h50;
	15'he78: q<=8'h0d;
	15'he79: q<=8'hbd;
	15'he7a: q<=8'hb9;
	15'he7b: q<=8'h02;
	15'he7c: q<=8'h38;
	15'he7d: q<=8'he9;
	15'he7e: q<=8'h01;
	15'he7f: q<=8'h29;
	15'he80: q<=8'h0f;
	15'he81: q<=8'h9d;
	15'he82: q<=8'hb9;
	15'he83: q<=8'h02;
	15'he84: q<=8'ha9;
	15'he85: q<=8'h87;
	15'he86: q<=8'h9d;
	15'he87: q<=8'hcc;
	15'he88: q<=8'h02;
	15'he89: q<=8'hb8;
	15'he8a: q<=8'h50;
	15'he8b: q<=8'h1e;
	15'he8c: q<=8'hbd;
	15'he8d: q<=8'h83;
	15'he8e: q<=8'h02;
	15'he8f: q<=8'h29;
	15'he90: q<=8'h40;
	15'he91: q<=8'hf0;
	15'he92: q<=8'h0b;
	15'he93: q<=8'hbd;
	15'he94: q<=8'hb9;
	15'he95: q<=8'h02;
	15'he96: q<=8'h18;
	15'he97: q<=8'h69;
	15'he98: q<=8'h01;
	15'he99: q<=8'h29;
	15'he9a: q<=8'h0f;
	15'he9b: q<=8'h9d;
	15'he9c: q<=8'hb9;
	15'he9d: q<=8'h02;
	15'he9e: q<=8'hbd;
	15'he9f: q<=8'h83;
	15'hea0: q<=8'h02;
	15'hea1: q<=8'hbc;
	15'hea2: q<=8'hb9;
	15'hea3: q<=8'h02;
	15'hea4: q<=8'h20;
	15'hea5: q<=8'hd7;
	15'hea6: q<=8'h9e;
	15'hea7: q<=8'h9d;
	15'hea8: q<=8'hcc;
	15'hea9: q<=8'h02;
	15'heaa: q<=8'h60;
	15'heab: q<=8'had;
	15'heac: q<=8'h11;
	15'head: q<=8'h01;
	15'heae: q<=8'hf0;
	15'heaf: q<=8'h26;
	15'heb0: q<=8'hbd;
	15'heb1: q<=8'h83;
	15'heb2: q<=8'h02;
	15'heb3: q<=8'h29;
	15'heb4: q<=8'h40;
	15'heb5: q<=8'hf0;
	15'heb6: q<=8'h12;
	15'heb7: q<=8'hbd;
	15'heb8: q<=8'hb9;
	15'heb9: q<=8'h02;
	15'heba: q<=8'hc9;
	15'hebb: q<=8'h0e;
	15'hebc: q<=8'h90;
	15'hebd: q<=8'h08;
	15'hebe: q<=8'hbd;
	15'hebf: q<=8'h83;
	15'hec0: q<=8'h02;
	15'hec1: q<=8'h29;
	15'hec2: q<=8'hbf;
	15'hec3: q<=8'h9d;
	15'hec4: q<=8'h83;
	15'hec5: q<=8'h02;
	15'hec6: q<=8'hb8;
	15'hec7: q<=8'h50;
	15'hec8: q<=8'h0d;
	15'hec9: q<=8'hbd;
	15'heca: q<=8'hb9;
	15'hecb: q<=8'h02;
	15'hecc: q<=8'hd0;
	15'hecd: q<=8'h08;
	15'hece: q<=8'hbd;
	15'hecf: q<=8'h83;
	15'hed0: q<=8'h02;
	15'hed1: q<=8'h09;
	15'hed2: q<=8'h40;
	15'hed3: q<=8'h9d;
	15'hed4: q<=8'h83;
	15'hed5: q<=8'h02;
	15'hed6: q<=8'h60;
	15'hed7: q<=8'h29;
	15'hed8: q<=8'h40;
	15'hed9: q<=8'hf0;
	15'heda: q<=8'h10;
	15'hedb: q<=8'h88;
	15'hedc: q<=8'h98;
	15'hedd: q<=8'h29;
	15'hede: q<=8'h0f;
	15'hedf: q<=8'ha8;
	15'hee0: q<=8'hb9;
	15'hee1: q<=8'hee;
	15'hee2: q<=8'h03;
	15'hee3: q<=8'h18;
	15'hee4: q<=8'h69;
	15'hee5: q<=8'h08;
	15'hee6: q<=8'h29;
	15'hee7: q<=8'h0f;
	15'hee8: q<=8'hb8;
	15'hee9: q<=8'h50;
	15'heea: q<=8'h03;
	15'heeb: q<=8'hb9;
	15'heec: q<=8'hee;
	15'heed: q<=8'h03;
	15'heee: q<=8'h09;
	15'heef: q<=8'h80;
	15'hef0: q<=8'h60;
	15'hef1: q<=8'ha0;
	15'hef2: q<=8'h04;
	15'hef3: q<=8'hbd;
	15'hef4: q<=8'h8a;
	15'hef5: q<=8'h02;
	15'hef6: q<=8'h30;
	15'hef7: q<=8'h4b;
	15'hef8: q<=8'hbd;
	15'hef9: q<=8'h9f;
	15'hefa: q<=8'h02;
	15'hefb: q<=8'h18;
	15'hefc: q<=8'h6d;
	15'hefd: q<=8'h64;
	15'hefe: q<=8'h01;
	15'heff: q<=8'h9d;
	15'hf00: q<=8'h9f;
	15'hf01: q<=8'h02;
	15'hf02: q<=8'hbd;
	15'hf03: q<=8'hdf;
	15'hf04: q<=8'h02;
	15'hf05: q<=8'h6d;
	15'hf06: q<=8'h69;
	15'hf07: q<=8'h01;
	15'hf08: q<=8'h9d;
	15'hf09: q<=8'hdf;
	15'hf0a: q<=8'h02;
	15'hf0b: q<=8'hcd;
	15'hf0c: q<=8'h02;
	15'hf0d: q<=8'h02;
	15'hf0e: q<=8'hb0;
	15'hf0f: q<=8'h09;
	15'hf10: q<=8'had;
	15'hf11: q<=8'h02;
	15'hf12: q<=8'h02;
	15'hf13: q<=8'h9d;
	15'hf14: q<=8'hdf;
	15'hf15: q<=8'h02;
	15'hf16: q<=8'hb8;
	15'hf17: q<=8'h50;
	15'hf18: q<=8'h11;
	15'hf19: q<=8'hac;
	15'hf1a: q<=8'hab;
	15'hf1b: q<=8'h03;
	15'hf1c: q<=8'hf0;
	15'hf1d: q<=8'h0b;
	15'hf1e: q<=8'ha4;
	15'hf1f: q<=8'h9f;
	15'hf20: q<=8'hc0;
	15'hf21: q<=8'h11;
	15'hf22: q<=8'hb0;
	15'hf23: q<=8'h02;
	15'hf24: q<=8'hc9;
	15'hf25: q<=8'h20;
	15'hf26: q<=8'hb8;
	15'hf27: q<=8'h50;
	15'hf28: q<=8'h01;
	15'hf29: q<=8'h60;
	15'hf2a: q<=8'hb0;
	15'hf2b: q<=8'h11;
	15'hf2c: q<=8'had;
	15'hf2d: q<=8'h59;
	15'hf2e: q<=8'h01;
	15'hf2f: q<=8'h10;
	15'hf30: q<=8'h06;
	15'hf31: q<=8'h20;
	15'hf32: q<=8'h81;
	15'hf33: q<=8'h9f;
	15'hf34: q<=8'hb8;
	15'hf35: q<=8'h50;
	15'hf36: q<=8'h03;
	15'hf37: q<=8'h20;
	15'hf38: q<=8'h8a;
	15'hf39: q<=8'h9f;
	15'hf3a: q<=8'hb8;
	15'hf3b: q<=8'h50;
	15'hf3c: q<=8'h03;
	15'hf3d: q<=8'h20;
	15'hf3e: q<=8'h5f;
	15'hf3f: q<=8'h9f;
	15'hf40: q<=8'hb8;
	15'hf41: q<=8'h50;
	15'hf42: q<=8'h1b;
	15'hf43: q<=8'h20;
	15'hf44: q<=8'h99;
	15'hf45: q<=8'h9c;
	15'hf46: q<=8'hc9;
	15'hf47: q<=8'h80;
	15'hf48: q<=8'h90;
	15'hf49: q<=8'h11;
	15'hf4a: q<=8'h2c;
	15'hf4b: q<=8'h59;
	15'hf4c: q<=8'h01;
	15'hf4d: q<=8'h50;
	15'hf4e: q<=8'h06;
	15'hf4f: q<=8'h20;
	15'hf50: q<=8'h81;
	15'hf51: q<=8'h9f;
	15'hf52: q<=8'hb8;
	15'hf53: q<=8'h50;
	15'hf54: q<=8'h03;
	15'hf55: q<=8'h20;
	15'hf56: q<=8'h8a;
	15'hf57: q<=8'h9f;
	15'hf58: q<=8'hb8;
	15'hf59: q<=8'h50;
	15'hf5a: q<=8'h03;
	15'hf5b: q<=8'h20;
	15'hf5c: q<=8'h5f;
	15'hf5d: q<=8'h9f;
	15'hf5e: q<=8'h60;
	15'hf5f: q<=8'hbd;
	15'hf60: q<=8'hdf;
	15'hf61: q<=8'h02;
	15'hf62: q<=8'h29;
	15'hf63: q<=8'h20;
	15'hf64: q<=8'hf0;
	15'hf65: q<=8'h1a;
	15'hf66: q<=8'had;
	15'hf67: q<=8'hda;
	15'hf68: q<=8'h60;
	15'hf69: q<=8'hcd;
	15'hf6a: q<=8'h5f;
	15'hf6b: q<=8'h01;
	15'hf6c: q<=8'h90;
	15'hf6d: q<=8'h12;
	15'hf6e: q<=8'h2c;
	15'hf6f: q<=8'h59;
	15'hf70: q<=8'h01;
	15'hf71: q<=8'h50;
	15'hf72: q<=8'h0a;
	15'hf73: q<=8'h8a;
	15'hf74: q<=8'h4a;
	15'hf75: q<=8'h90;
	15'hf76: q<=8'h13;
	15'hf77: q<=8'h20;
	15'hf78: q<=8'h81;
	15'hf79: q<=8'h9f;
	15'hf7a: q<=8'hb8;
	15'hf7b: q<=8'h50;
	15'hf7c: q<=8'h03;
	15'hf7d: q<=8'h20;
	15'hf7e: q<=8'h8a;
	15'hf7f: q<=8'h9f;
	15'hf80: q<=8'h60;
	15'hf81: q<=8'h20;
	15'hf82: q<=8'h67;
	15'hf83: q<=8'h9d;
	15'hf84: q<=8'h20;
	15'hf85: q<=8'h4f;
	15'hf86: q<=8'h9c;
	15'hf87: q<=8'h4c;
	15'hf88: q<=8'h99;
	15'hf89: q<=8'h9f;
	15'hf8a: q<=8'hbd;
	15'hf8b: q<=8'h83;
	15'hf8c: q<=8'h02;
	15'hf8d: q<=8'h29;
	15'hf8e: q<=8'hbf;
	15'hf8f: q<=8'h2c;
	15'hf90: q<=8'hca;
	15'hf91: q<=8'h60;
	15'hf92: q<=8'h50;
	15'hf93: q<=8'h02;
	15'hf94: q<=8'h09;
	15'hf95: q<=8'h40;
	15'hf96: q<=8'h9d;
	15'hf97: q<=8'h83;
	15'hf98: q<=8'h02;
	15'hf99: q<=8'had;
	15'hf9a: q<=8'h11;
	15'hf9b: q<=8'h01;
	15'hf9c: q<=8'hf0;
	15'hf9d: q<=8'h1e;
	15'hf9e: q<=8'hbd;
	15'hf9f: q<=8'h83;
	15'hfa0: q<=8'h02;
	15'hfa1: q<=8'h29;
	15'hfa2: q<=8'h40;
	15'hfa3: q<=8'hd0;
	15'hfa4: q<=8'h0a;
	15'hfa5: q<=8'hbd;
	15'hfa6: q<=8'hb9;
	15'hfa7: q<=8'h02;
	15'hfa8: q<=8'hc9;
	15'hfa9: q<=8'h0f;
	15'hfaa: q<=8'hb0;
	15'hfab: q<=8'h08;
	15'hfac: q<=8'hb8;
	15'hfad: q<=8'h50;
	15'hfae: q<=8'h0d;
	15'hfaf: q<=8'hbd;
	15'hfb0: q<=8'hb9;
	15'hfb1: q<=8'h02;
	15'hfb2: q<=8'hd0;
	15'hfb3: q<=8'h08;
	15'hfb4: q<=8'hbd;
	15'hfb5: q<=8'h83;
	15'hfb6: q<=8'h02;
	15'hfb7: q<=8'h49;
	15'hfb8: q<=8'h40;
	15'hfb9: q<=8'h9d;
	15'hfba: q<=8'h83;
	15'hfbb: q<=8'h02;
	15'hfbc: q<=8'ha9;
	15'hfbd: q<=8'h66;
	15'hfbe: q<=8'h8d;
	15'hfbf: q<=8'h0b;
	15'hfc0: q<=8'h01;
	15'hfc1: q<=8'h4c;
	15'hfc2: q<=8'h5f;
	15'hfc3: q<=8'h9e;
	15'hfc4: q<=8'ha9;
	15'hfc5: q<=8'h01;
	15'hfc6: q<=8'h8d;
	15'hfc7: q<=8'h0c;
	15'hfc8: q<=8'h01;
	15'hfc9: q<=8'hbc;
	15'hfca: q<=8'hb9;
	15'hfcb: q<=8'h02;
	15'hfcc: q<=8'hb9;
	15'hfcd: q<=8'hac;
	15'hfce: q<=8'h03;
	15'hfcf: q<=8'hd0;
	15'hfd0: q<=8'h05;
	15'hfd1: q<=8'ha9;
	15'hfd2: q<=8'hf1;
	15'hfd3: q<=8'h99;
	15'hfd4: q<=8'hac;
	15'hfd5: q<=8'h03;
	15'hfd6: q<=8'hbd;
	15'hfd7: q<=8'hdf;
	15'hfd8: q<=8'h02;
	15'hfd9: q<=8'hd9;
	15'hfda: q<=8'hac;
	15'hfdb: q<=8'h03;
	15'hfdc: q<=8'hb0;
	15'hfdd: q<=8'h08;
	15'hfde: q<=8'h99;
	15'hfdf: q<=8'hac;
	15'hfe0: q<=8'h03;
	15'hfe1: q<=8'ha9;
	15'hfe2: q<=8'h80;
	15'hfe3: q<=8'h99;
	15'hfe4: q<=8'h9a;
	15'hfe5: q<=8'h03;
	15'hfe6: q<=8'hbd;
	15'hfe7: q<=8'hdf;
	15'hfe8: q<=8'h02;
	15'hfe9: q<=8'hc9;
	15'hfea: q<=8'h20;
	15'hfeb: q<=8'hb0;
	15'hfec: q<=8'h10;
	15'hfed: q<=8'hbd;
	15'hfee: q<=8'h8a;
	15'hfef: q<=8'h02;
	15'hff0: q<=8'h09;
	15'hff1: q<=8'h80;
	15'hff2: q<=8'h9d;
	15'hff3: q<=8'h8a;
	15'hff4: q<=8'h02;
	15'hff5: q<=8'ha9;
	15'hff6: q<=8'h20;
	15'hff7: q<=8'h9d;
	15'hff8: q<=8'hdf;
	15'hff9: q<=8'h02;
	15'hffa: q<=8'hb8;
	15'hffb: q<=8'h50;
	15'hffc: q<=8'h2a;
	15'hffd: q<=8'hc9;
	15'hffe: q<=8'hf2;
	15'hfff: q<=8'h90;
	15'h1000: q<=8'h26;
	15'h1001: q<=8'h20;
	15'h1002: q<=8'h28;
	15'h1003: q<=8'ha0;
	15'h1004: q<=8'ha9;
	15'h1005: q<=8'hf0;
	15'h1006: q<=8'h9d;
	15'h1007: q<=8'hdf;
	15'h1008: q<=8'h02;
	15'h1009: q<=8'had;
	15'h100a: q<=8'hab;
	15'h100b: q<=8'h03;
	15'h100c: q<=8'hd0;
	15'h100d: q<=8'h19;
	15'h100e: q<=8'hbd;
	15'h100f: q<=8'h8a;
	15'h1010: q<=8'h02;
	15'h1011: q<=8'h29;
	15'h1012: q<=8'hfc;
	15'h1013: q<=8'h09;
	15'h1014: q<=8'h01;
	15'h1015: q<=8'h9d;
	15'h1016: q<=8'h8a;
	15'h1017: q<=8'h02;
	15'h1018: q<=8'hbd;
	15'h1019: q<=8'h83;
	15'h101a: q<=8'h02;
	15'h101b: q<=8'h29;
	15'h101c: q<=8'hf8;
	15'h101d: q<=8'h09;
	15'h101e: q<=8'h02;
	15'h101f: q<=8'h9d;
	15'h1020: q<=8'h83;
	15'h1021: q<=8'h02;
	15'h1022: q<=8'ha9;
	15'h1023: q<=8'h00;
	15'h1024: q<=8'h8d;
	15'h1025: q<=8'h0c;
	15'h1026: q<=8'h01;
	15'h1027: q<=8'h60;
	15'h1028: q<=8'ha9;
	15'h1029: q<=8'h00;
	15'h102a: q<=8'h85;
	15'h102b: q<=8'h2d;
	15'h102c: q<=8'ha9;
	15'h102d: q<=8'h0f;
	15'h102e: q<=8'h8d;
	15'h102f: q<=8'h40;
	15'h1030: q<=8'h01;
	15'h1031: q<=8'had;
	15'h1032: q<=8'hda;
	15'h1033: q<=8'h60;
	15'h1034: q<=8'h29;
	15'h1035: q<=8'h0f;
	15'h1036: q<=8'ha8;
	15'h1037: q<=8'hc0;
	15'h1038: q<=8'h0f;
	15'h1039: q<=8'hd0;
	15'h103a: q<=8'h05;
	15'h103b: q<=8'had;
	15'h103c: q<=8'h11;
	15'h103d: q<=8'h01;
	15'h103e: q<=8'hd0;
	15'h103f: q<=8'h0f;
	15'h1040: q<=8'hb9;
	15'h1041: q<=8'hac;
	15'h1042: q<=8'h03;
	15'h1043: q<=8'hd0;
	15'h1044: q<=8'h02;
	15'h1045: q<=8'ha9;
	15'h1046: q<=8'hff;
	15'h1047: q<=8'hc5;
	15'h1048: q<=8'h2d;
	15'h1049: q<=8'h90;
	15'h104a: q<=8'h04;
	15'h104b: q<=8'h85;
	15'h104c: q<=8'h2d;
	15'h104d: q<=8'h84;
	15'h104e: q<=8'h29;
	15'h104f: q<=8'h88;
	15'h1050: q<=8'h10;
	15'h1051: q<=8'h02;
	15'h1052: q<=8'ha0;
	15'h1053: q<=8'h0f;
	15'h1054: q<=8'hce;
	15'h1055: q<=8'h40;
	15'h1056: q<=8'h01;
	15'h1057: q<=8'h10;
	15'h1058: q<=8'hde;
	15'h1059: q<=8'ha5;
	15'h105a: q<=8'h29;
	15'h105b: q<=8'h9d;
	15'h105c: q<=8'hb9;
	15'h105d: q<=8'h02;
	15'h105e: q<=8'h18;
	15'h105f: q<=8'h69;
	15'h1060: q<=8'h01;
	15'h1061: q<=8'h29;
	15'h1062: q<=8'h0f;
	15'h1063: q<=8'h9d;
	15'h1064: q<=8'hcc;
	15'h1065: q<=8'h02;
	15'h1066: q<=8'hbd;
	15'h1067: q<=8'h8a;
	15'h1068: q<=8'h02;
	15'h1069: q<=8'h29;
	15'h106a: q<=8'h7f;
	15'h106b: q<=8'h9d;
	15'h106c: q<=8'h8a;
	15'h106d: q<=8'h02;
	15'h106e: q<=8'h60;
	15'h106f: q<=8'hb9;
	15'h1070: q<=8'hdf;
	15'h1071: q<=8'h02;
	15'h1072: q<=8'h85;
	15'h1073: q<=8'h29;
	15'h1074: q<=8'hcd;
	15'h1075: q<=8'h02;
	15'h1076: q<=8'h02;
	15'h1077: q<=8'hd0;
	15'h1078: q<=8'h0f;
	15'h1079: q<=8'hb9;
	15'h107a: q<=8'h83;
	15'h107b: q<=8'h02;
	15'h107c: q<=8'h29;
	15'h107d: q<=8'h07;
	15'h107e: q<=8'hc9;
	15'h107f: q<=8'h04;
	15'h1080: q<=8'hf0;
	15'h1081: q<=8'h06;
	15'h1082: q<=8'hce;
	15'h1083: q<=8'h09;
	15'h1084: q<=8'h01;
	15'h1085: q<=8'hb8;
	15'h1086: q<=8'h50;
	15'h1087: q<=8'h03;
	15'h1088: q<=8'hce;
	15'h1089: q<=8'h08;
	15'h108a: q<=8'h01;
	15'h108b: q<=8'ha9;
	15'h108c: q<=8'h00;
	15'h108d: q<=8'h99;
	15'h108e: q<=8'hdf;
	15'h108f: q<=8'h02;
	15'h1090: q<=8'hb9;
	15'h1091: q<=8'h83;
	15'h1092: q<=8'h02;
	15'h1093: q<=8'h29;
	15'h1094: q<=8'h07;
	15'h1095: q<=8'h86;
	15'h1096: q<=8'h35;
	15'h1097: q<=8'haa;
	15'h1098: q<=8'hde;
	15'h1099: q<=8'h42;
	15'h109a: q<=8'h01;
	15'h109b: q<=8'ha6;
	15'h109c: q<=8'h35;
	15'h109d: q<=8'hb9;
	15'h109e: q<=8'h8a;
	15'h109f: q<=8'h02;
	15'h10a0: q<=8'h29;
	15'h10a1: q<=8'h03;
	15'h10a2: q<=8'hf0;
	15'h10a3: q<=8'h52;
	15'h10a4: q<=8'h38;
	15'h10a5: q<=8'he9;
	15'h10a6: q<=8'h01;
	15'h10a7: q<=8'hc9;
	15'h10a8: q<=8'h02;
	15'h10a9: q<=8'hd0;
	15'h10aa: q<=8'h02;
	15'h10ab: q<=8'ha9;
	15'h10ac: q<=8'h04;
	15'h10ad: q<=8'h85;
	15'h10ae: q<=8'h2b;
	15'h10af: q<=8'hb9;
	15'h10b0: q<=8'hb9;
	15'h10b1: q<=8'h02;
	15'h10b2: q<=8'h38;
	15'h10b3: q<=8'he9;
	15'h10b4: q<=8'h01;
	15'h10b5: q<=8'h29;
	15'h10b6: q<=8'h0f;
	15'h10b7: q<=8'hc9;
	15'h10b8: q<=8'h0f;
	15'h10b9: q<=8'h90;
	15'h10ba: q<=8'h07;
	15'h10bb: q<=8'h2c;
	15'h10bc: q<=8'h11;
	15'h10bd: q<=8'h01;
	15'h10be: q<=8'h10;
	15'h10bf: q<=8'h02;
	15'h10c0: q<=8'ha9;
	15'h10c1: q<=8'h00;
	15'h10c2: q<=8'h85;
	15'h10c3: q<=8'h2a;
	15'h10c4: q<=8'h20;
	15'h10c5: q<=8'h07;
	15'h10c6: q<=8'h9b;
	15'h10c7: q<=8'ha5;
	15'h10c8: q<=8'h2d;
	15'h10c9: q<=8'h8d;
	15'h10ca: q<=8'h0b;
	15'h10cb: q<=8'h01;
	15'h10cc: q<=8'hce;
	15'h10cd: q<=8'h0b;
	15'h10ce: q<=8'h01;
	15'h10cf: q<=8'ha9;
	15'h10d0: q<=8'h00;
	15'h10d1: q<=8'h8d;
	15'h10d2: q<=8'h0a;
	15'h10d3: q<=8'h01;
	15'h10d4: q<=8'h20;
	15'h10d5: q<=8'h4d;
	15'h10d6: q<=8'h99;
	15'h10d7: q<=8'hf0;
	15'h10d8: q<=8'h1d;
	15'h10d9: q<=8'ha5;
	15'h10da: q<=8'h2a;
	15'h10db: q<=8'h18;
	15'h10dc: q<=8'h69;
	15'h10dd: q<=8'h02;
	15'h10de: q<=8'h29;
	15'h10df: q<=8'h0f;
	15'h10e0: q<=8'hc9;
	15'h10e1: q<=8'h0f;
	15'h10e2: q<=8'hd0;
	15'h10e3: q<=8'h07;
	15'h10e4: q<=8'h2c;
	15'h10e5: q<=8'h11;
	15'h10e6: q<=8'h01;
	15'h10e7: q<=8'h10;
	15'h10e8: q<=8'h02;
	15'h10e9: q<=8'ha9;
	15'h10ea: q<=8'h0e;
	15'h10eb: q<=8'h85;
	15'h10ec: q<=8'h2a;
	15'h10ed: q<=8'ha5;
	15'h10ee: q<=8'h2b;
	15'h10ef: q<=8'h09;
	15'h10f0: q<=8'h40;
	15'h10f1: q<=8'h85;
	15'h10f2: q<=8'h2b;
	15'h10f3: q<=8'h20;
	15'h10f4: q<=8'h4d;
	15'h10f5: q<=8'h99;
	15'h10f6: q<=8'h60;
	15'h10f7: q<=8'h0c;
	15'h10f8: q<=8'h0e;
	15'h10f9: q<=8'h1a;
	15'h10fa: q<=8'h06;
	15'h10fb: q<=8'h00;
	15'h10fc: q<=8'h06;
	15'h10fd: q<=8'hff;
	15'h10fe: q<=8'h0c;
	15'h10ff: q<=8'h00;
	15'h1100: q<=8'h06;
	15'h1101: q<=8'h06;
	15'h1102: q<=8'h02;
	15'h1103: q<=8'h08;
	15'h1104: q<=8'h0c;
	15'h1105: q<=8'h00;
	15'h1106: q<=8'h08;
	15'h1107: q<=8'h0c;
	15'h1108: q<=8'h12;
	15'h1109: q<=8'h00;
	15'h110a: q<=8'h14;
	15'h110b: q<=8'h04;
	15'h110c: q<=8'h06;
	15'h110d: q<=8'h11;
	15'h110e: q<=8'h06;
	15'h110f: q<=8'h0a;
	15'h1110: q<=8'h0c;
	15'h1111: q<=8'h00;
	15'h1112: q<=8'h12;
	15'h1113: q<=8'h00;
	15'h1114: q<=8'h14;
	15'h1115: q<=8'h0c;
	15'h1116: q<=8'h04;
	15'h1117: q<=8'h06;
	15'h1118: q<=8'h1b;
	15'h1119: q<=8'h06;
	15'h111a: q<=8'h18;
	15'h111b: q<=8'h0c;
	15'h111c: q<=8'h00;
	15'h111d: q<=8'h02;
	15'h111e: q<=8'h02;
	15'h111f: q<=8'h12;
	15'h1120: q<=8'h00;
	15'h1121: q<=8'h14;
	15'h1122: q<=8'h0c;
	15'h1123: q<=8'h04;
	15'h1124: q<=8'h06;
	15'h1125: q<=8'h28;
	15'h1126: q<=8'h00;
	15'h1127: q<=8'h08;
	15'h1128: q<=8'h27;
	15'h1129: q<=8'h16;
	15'h112a: q<=8'h02;
	15'h112b: q<=8'h03;
	15'h112c: q<=8'h12;
	15'h112d: q<=8'h00;
	15'h112e: q<=8'h14;
	15'h112f: q<=8'h0c;
	15'h1130: q<=8'h04;
	15'h1131: q<=8'h06;
	15'h1132: q<=8'h35;
	15'h1133: q<=8'h00;
	15'h1134: q<=8'h08;
	15'h1135: q<=8'h34;
	15'h1136: q<=8'h16;
	15'h1137: q<=8'h06;
	15'h1138: q<=8'h23;
	15'h1139: q<=8'h02;
	15'h113a: q<=8'h04;
	15'h113b: q<=8'h18;
	15'h113c: q<=8'h00;
	15'h113d: q<=8'h08;
	15'h113e: q<=8'h43;
	15'h113f: q<=8'h12;
	15'h1140: q<=8'h00;
	15'h1141: q<=8'h10;
	15'h1142: q<=8'hb3;
	15'h1143: q<=8'h14;
	15'h1144: q<=8'h1a;
	15'h1145: q<=8'h41;
	15'h1146: q<=8'h08;
	15'h1147: q<=8'h4b;
	15'h1148: q<=8'h06;
	15'h1149: q<=8'h48;
	15'h114a: q<=8'h00;
	15'h114b: q<=8'h0c;
	15'h114c: q<=8'h1c;
	15'h114d: q<=8'h1a;
	15'h114e: q<=8'h52;
	15'h114f: q<=8'h12;
	15'h1150: q<=8'h00;
	15'h1151: q<=8'h0c;
	15'h1152: q<=8'h14;
	15'h1153: q<=8'h1a;
	15'h1154: q<=8'h52;
	15'h1155: q<=8'h00;
	15'h1156: q<=8'h06;
	15'h1157: q<=8'h5a;
	15'h1158: q<=8'h1e;
	15'h1159: q<=8'h20;
	15'h115a: q<=8'h00;
	15'h115b: q<=8'h06;
	15'h115c: q<=8'h60;
	15'h115d: q<=8'h00;
	15'h115e: q<=8'h02;
	15'h115f: q<=8'h03;
	15'h1160: q<=8'h20;
	15'h1161: q<=8'h00;
	15'h1162: q<=8'h08;
	15'h1163: q<=8'h68;
	15'h1164: q<=8'h14;
	15'h1165: q<=8'h1a;
	15'h1166: q<=8'h60;
	15'h1167: q<=8'h06;
	15'h1168: q<=8'h65;
	15'h1169: q<=8'h10;
	15'h116a: q<=8'hb2;
	15'h116b: q<=8'h22;
	15'h116c: q<=8'h00;
	15'h116d: q<=8'h08;
	15'h116e: q<=8'h73;
	15'h116f: q<=8'h26;
	15'h1170: q<=8'h1a;
	15'h1171: q<=8'h7e;
	15'h1172: q<=8'h22;
	15'h1173: q<=8'h00;
	15'h1174: q<=8'h06;
	15'h1175: q<=8'h77;
	15'h1176: q<=8'h24;
	15'h1177: q<=8'h12;
	15'h1178: q<=8'h00;
	15'h1179: q<=8'h14;
	15'h117a: q<=8'h1a;
	15'h117b: q<=8'h71;
	15'h117c: q<=8'h06;
	15'h117d: q<=8'h80;
	15'h117e: q<=8'h24;
	15'h117f: q<=8'h16;
	15'h1180: q<=8'h12;
	15'h1181: q<=8'h00;
	15'h1182: q<=8'h0c;
	15'h1183: q<=8'h14;
	15'h1184: q<=8'h04;
	15'h1185: q<=8'h06;
	15'h1186: q<=8'h89;
	15'h1187: q<=8'h02;
	15'h1188: q<=8'h04;
	15'h1189: q<=8'h00;
	15'h118a: q<=8'h0c;
	15'h118b: q<=8'h08;
	15'h118c: q<=8'h91;
	15'h118d: q<=8'h06;
	15'h118e: q<=8'h86;
	15'h118f: q<=8'ha2;
	15'h1190: q<=8'h0b;
	15'h1191: q<=8'h86;
	15'h1192: q<=8'h37;
	15'h1193: q<=8'ha6;
	15'h1194: q<=8'h37;
	15'h1195: q<=8'hbd;
	15'h1196: q<=8'hd3;
	15'h1197: q<=8'h02;
	15'h1198: q<=8'hf0;
	15'h1199: q<=8'h45;
	15'h119a: q<=8'he0;
	15'h119b: q<=8'h08;
	15'h119c: q<=8'hb0;
	15'h119d: q<=8'h22;
	15'h119e: q<=8'h69;
	15'h119f: q<=8'h09;
	15'h11a0: q<=8'hbc;
	15'h11a1: q<=8'hf2;
	15'h11a2: q<=8'h02;
	15'h11a3: q<=8'hf0;
	15'h11a4: q<=8'h03;
	15'h11a5: q<=8'h38;
	15'h11a6: q<=8'he9;
	15'h11a7: q<=8'h04;
	15'h11a8: q<=8'h9d;
	15'h11a9: q<=8'hd3;
	15'h11aa: q<=8'h02;
	15'h11ab: q<=8'h20;
	15'h11ac: q<=8'hfa;
	15'h11ad: q<=8'ha1;
	15'h11ae: q<=8'hbd;
	15'h11af: q<=8'hd3;
	15'h11b0: q<=8'h02;
	15'h11b1: q<=8'hc9;
	15'h11b2: q<=8'hf0;
	15'h11b3: q<=8'h90;
	15'h11b4: q<=8'h08;
	15'h11b5: q<=8'hce;
	15'h11b6: q<=8'h35;
	15'h11b7: q<=8'h01;
	15'h11b8: q<=8'ha9;
	15'h11b9: q<=8'h00;
	15'h11ba: q<=8'h9d;
	15'h11bb: q<=8'hd3;
	15'h11bc: q<=8'h02;
	15'h11bd: q<=8'hb8;
	15'h11be: q<=8'h50;
	15'h11bf: q<=8'h1f;
	15'h11c0: q<=8'hbd;
	15'h11c1: q<=8'he6;
	15'h11c2: q<=8'h02;
	15'h11c3: q<=8'h18;
	15'h11c4: q<=8'h6d;
	15'h11c5: q<=8'h20;
	15'h11c6: q<=8'h01;
	15'h11c7: q<=8'h9d;
	15'h11c8: q<=8'he6;
	15'h11c9: q<=8'h02;
	15'h11ca: q<=8'hbd;
	15'h11cb: q<=8'hd3;
	15'h11cc: q<=8'h02;
	15'h11cd: q<=8'h6d;
	15'h11ce: q<=8'h18;
	15'h11cf: q<=8'h01;
	15'h11d0: q<=8'hcd;
	15'h11d1: q<=8'h02;
	15'h11d2: q<=8'h02;
	15'h11d3: q<=8'hb0;
	15'h11d4: q<=8'h07;
	15'h11d5: q<=8'hc6;
	15'h11d6: q<=8'ha6;
	15'h11d7: q<=8'h20;
	15'h11d8: q<=8'he4;
	15'h11d9: q<=8'ha1;
	15'h11da: q<=8'ha9;
	15'h11db: q<=8'h00;
	15'h11dc: q<=8'h9d;
	15'h11dd: q<=8'hd3;
	15'h11de: q<=8'h02;
	15'h11df: q<=8'hc6;
	15'h11e0: q<=8'h37;
	15'h11e1: q<=8'h10;
	15'h11e2: q<=8'hb0;
	15'h11e3: q<=8'h60;
	15'h11e4: q<=8'had;
	15'h11e5: q<=8'h00;
	15'h11e6: q<=8'h02;
	15'h11e7: q<=8'hdd;
	15'h11e8: q<=8'had;
	15'h11e9: q<=8'h02;
	15'h11ea: q<=8'hd0;
	15'h11eb: q<=8'h0d;
	15'h11ec: q<=8'had;
	15'h11ed: q<=8'h01;
	15'h11ee: q<=8'h02;
	15'h11ef: q<=8'h30;
	15'h11f0: q<=8'h08;
	15'h11f1: q<=8'h20;
	15'h11f2: q<=8'h4b;
	15'h11f3: q<=8'ha3;
	15'h11f4: q<=8'ha9;
	15'h11f5: q<=8'h81;
	15'h11f6: q<=8'h8d;
	15'h11f7: q<=8'h01;
	15'h11f8: q<=8'h02;
	15'h11f9: q<=8'h60;
	15'h11fa: q<=8'hbc;
	15'h11fb: q<=8'had;
	15'h11fc: q<=8'h02;
	15'h11fd: q<=8'hb9;
	15'h11fe: q<=8'hac;
	15'h11ff: q<=8'h03;
	15'h1200: q<=8'hf0;
	15'h1201: q<=8'h3c;
	15'h1202: q<=8'hbd;
	15'h1203: q<=8'hd3;
	15'h1204: q<=8'h02;
	15'h1205: q<=8'hd9;
	15'h1206: q<=8'hac;
	15'h1207: q<=8'h03;
	15'h1208: q<=8'h90;
	15'h1209: q<=8'h25;
	15'h120a: q<=8'hc9;
	15'h120b: q<=8'hf0;
	15'h120c: q<=8'h90;
	15'h120d: q<=8'h02;
	15'h120e: q<=8'ha9;
	15'h120f: q<=8'h00;
	15'h1210: q<=8'h99;
	15'h1211: q<=8'hac;
	15'h1212: q<=8'h03;
	15'h1213: q<=8'hfe;
	15'h1214: q<=8'hf2;
	15'h1215: q<=8'h02;
	15'h1216: q<=8'ha9;
	15'h1217: q<=8'hc0;
	15'h1218: q<=8'h99;
	15'h1219: q<=8'h9a;
	15'h121a: q<=8'h03;
	15'h121b: q<=8'h20;
	15'h121c: q<=8'hf6;
	15'h121d: q<=8'hcc;
	15'h121e: q<=8'ha2;
	15'h121f: q<=8'hff;
	15'h1220: q<=8'ha9;
	15'h1221: q<=8'h00;
	15'h1222: q<=8'h85;
	15'h1223: q<=8'h2a;
	15'h1224: q<=8'h85;
	15'h1225: q<=8'h2b;
	15'h1226: q<=8'ha9;
	15'h1227: q<=8'h01;
	15'h1228: q<=8'h85;
	15'h1229: q<=8'h29;
	15'h122a: q<=8'h20;
	15'h122b: q<=8'h6c;
	15'h122c: q<=8'hca;
	15'h122d: q<=8'ha6;
	15'h122e: q<=8'h37;
	15'h122f: q<=8'hbd;
	15'h1230: q<=8'hf2;
	15'h1231: q<=8'h02;
	15'h1232: q<=8'hc9;
	15'h1233: q<=8'h02;
	15'h1234: q<=8'h90;
	15'h1235: q<=8'h08;
	15'h1236: q<=8'ha9;
	15'h1237: q<=8'h00;
	15'h1238: q<=8'h9d;
	15'h1239: q<=8'hd3;
	15'h123a: q<=8'h02;
	15'h123b: q<=8'hce;
	15'h123c: q<=8'h35;
	15'h123d: q<=8'h01;
	15'h123e: q<=8'h60;
	15'h123f: q<=8'had;
	15'h1240: q<=8'h01;
	15'h1241: q<=8'h02;
	15'h1242: q<=8'h30;
	15'h1243: q<=8'h61;
	15'h1244: q<=8'ha5;
	15'h1245: q<=8'h05;
	15'h1246: q<=8'h30;
	15'h1247: q<=8'h28;
	15'h1248: q<=8'had;
	15'h1249: q<=8'h06;
	15'h124a: q<=8'h01;
	15'h124b: q<=8'h85;
	15'h124c: q<=8'h29;
	15'h124d: q<=8'ha2;
	15'h124e: q<=8'h0a;
	15'h124f: q<=8'hbd;
	15'h1250: q<=8'hdb;
	15'h1251: q<=8'h02;
	15'h1252: q<=8'hf0;
	15'h1253: q<=8'h14;
	15'h1254: q<=8'hbd;
	15'h1255: q<=8'hb5;
	15'h1256: q<=8'h02;
	15'h1257: q<=8'h38;
	15'h1258: q<=8'hed;
	15'h1259: q<=8'h00;
	15'h125a: q<=8'h02;
	15'h125b: q<=8'h10;
	15'h125c: q<=8'h05;
	15'h125d: q<=8'h49;
	15'h125e: q<=8'hff;
	15'h125f: q<=8'h18;
	15'h1260: q<=8'h69;
	15'h1261: q<=8'h01;
	15'h1262: q<=8'hc9;
	15'h1263: q<=8'h02;
	15'h1264: q<=8'hb0;
	15'h1265: q<=8'h02;
	15'h1266: q<=8'he6;
	15'h1267: q<=8'h29;
	15'h1268: q<=8'hca;
	15'h1269: q<=8'h10;
	15'h126a: q<=8'he4;
	15'h126b: q<=8'ha5;
	15'h126c: q<=8'h29;
	15'h126d: q<=8'hb8;
	15'h126e: q<=8'h50;
	15'h126f: q<=8'h04;
	15'h1270: q<=8'ha5;
	15'h1271: q<=8'h4d;
	15'h1272: q<=8'h29;
	15'h1273: q<=8'h10;
	15'h1274: q<=8'hf0;
	15'h1275: q<=8'h2f;
	15'h1276: q<=8'ha2;
	15'h1277: q<=8'h07;
	15'h1278: q<=8'hbd;
	15'h1279: q<=8'hd3;
	15'h127a: q<=8'h02;
	15'h127b: q<=8'hd0;
	15'h127c: q<=8'h25;
	15'h127d: q<=8'hee;
	15'h127e: q<=8'h35;
	15'h127f: q<=8'h01;
	15'h1280: q<=8'had;
	15'h1281: q<=8'h02;
	15'h1282: q<=8'h02;
	15'h1283: q<=8'h9d;
	15'h1284: q<=8'hd3;
	15'h1285: q<=8'h02;
	15'h1286: q<=8'had;
	15'h1287: q<=8'h00;
	15'h1288: q<=8'h02;
	15'h1289: q<=8'h9d;
	15'h128a: q<=8'had;
	15'h128b: q<=8'h02;
	15'h128c: q<=8'had;
	15'h128d: q<=8'h01;
	15'h128e: q<=8'h02;
	15'h128f: q<=8'h9d;
	15'h1290: q<=8'hc0;
	15'h1291: q<=8'h02;
	15'h1292: q<=8'ha9;
	15'h1293: q<=8'h00;
	15'h1294: q<=8'h9d;
	15'h1295: q<=8'hf2;
	15'h1296: q<=8'h02;
	15'h1297: q<=8'h20;
	15'h1298: q<=8'hea;
	15'h1299: q<=8'hcc;
	15'h129a: q<=8'had;
	15'h129b: q<=8'h02;
	15'h129c: q<=8'h02;
	15'h129d: q<=8'h20;
	15'h129e: q<=8'h63;
	15'h129f: q<=8'ha4;
	15'h12a0: q<=8'ha2;
	15'h12a1: q<=8'h00;
	15'h12a2: q<=8'hca;
	15'h12a3: q<=8'h10;
	15'h12a4: q<=8'hd3;
	15'h12a5: q<=8'h60;
	15'h12a6: q<=8'had;
	15'h12a7: q<=8'h01;
	15'h12a8: q<=8'h02;
	15'h12a9: q<=8'h30;
	15'h12aa: q<=8'h58;
	15'h12ab: q<=8'ha2;
	15'h12ac: q<=8'h06;
	15'h12ad: q<=8'hbd;
	15'h12ae: q<=8'hdf;
	15'h12af: q<=8'h02;
	15'h12b0: q<=8'hf0;
	15'h12b1: q<=8'h4e;
	15'h12b2: q<=8'hc9;
	15'h12b3: q<=8'h30;
	15'h12b4: q<=8'h90;
	15'h12b5: q<=8'h4a;
	15'h12b6: q<=8'hbd;
	15'h12b7: q<=8'h8a;
	15'h12b8: q<=8'h02;
	15'h12b9: q<=8'h29;
	15'h12ba: q<=8'h40;
	15'h12bb: q<=8'hf0;
	15'h12bc: q<=8'h43;
	15'h12bd: q<=8'hde;
	15'h12be: q<=8'ha6;
	15'h12bf: q<=8'h02;
	15'h12c0: q<=8'h10;
	15'h12c1: q<=8'h3e;
	15'h12c2: q<=8'hfe;
	15'h12c3: q<=8'ha6;
	15'h12c4: q<=8'h02;
	15'h12c5: q<=8'hbd;
	15'h12c6: q<=8'h83;
	15'h12c7: q<=8'h02;
	15'h12c8: q<=8'h29;
	15'h12c9: q<=8'h80;
	15'h12ca: q<=8'hd0;
	15'h12cb: q<=8'h34;
	15'h12cc: q<=8'had;
	15'h12cd: q<=8'hca;
	15'h12ce: q<=8'h60;
	15'h12cf: q<=8'ha4;
	15'h12d0: q<=8'ha6;
	15'h12d1: q<=8'hd9;
	15'h12d2: q<=8'h04;
	15'h12d3: q<=8'ha3;
	15'h12d4: q<=8'h90;
	15'h12d5: q<=8'h2a;
	15'h12d6: q<=8'hac;
	15'h12d7: q<=8'h1a;
	15'h12d8: q<=8'h01;
	15'h12d9: q<=8'hb9;
	15'h12da: q<=8'hdb;
	15'h12db: q<=8'h02;
	15'h12dc: q<=8'hd0;
	15'h12dd: q<=8'h1f;
	15'h12de: q<=8'hbd;
	15'h12df: q<=8'hdf;
	15'h12e0: q<=8'h02;
	15'h12e1: q<=8'h99;
	15'h12e2: q<=8'hdb;
	15'h12e3: q<=8'h02;
	15'h12e4: q<=8'hbd;
	15'h12e5: q<=8'hb9;
	15'h12e6: q<=8'h02;
	15'h12e7: q<=8'h99;
	15'h12e8: q<=8'hb5;
	15'h12e9: q<=8'h02;
	15'h12ea: q<=8'hbd;
	15'h12eb: q<=8'hcc;
	15'h12ec: q<=8'h02;
	15'h12ed: q<=8'h99;
	15'h12ee: q<=8'hc8;
	15'h12ef: q<=8'h02;
	15'h12f0: q<=8'had;
	15'h12f1: q<=8'h19;
	15'h12f2: q<=8'h01;
	15'h12f3: q<=8'h9d;
	15'h12f4: q<=8'ha6;
	15'h12f5: q<=8'h02;
	15'h12f6: q<=8'h20;
	15'h12f7: q<=8'hbd;
	15'h12f8: q<=8'hcc;
	15'h12f9: q<=8'he6;
	15'h12fa: q<=8'ha6;
	15'h12fb: q<=8'ha0;
	15'h12fc: q<=8'h00;
	15'h12fd: q<=8'h88;
	15'h12fe: q<=8'h10;
	15'h12ff: q<=8'hd9;
	15'h1300: q<=8'hca;
	15'h1301: q<=8'h10;
	15'h1302: q<=8'haa;
	15'h1303: q<=8'h60;
	15'h1304: q<=8'h00;
	15'h1305: q<=8'he0;
	15'h1306: q<=8'hf0;
	15'h1307: q<=8'hfa;
	15'h1308: q<=8'hff;
	15'h1309: q<=8'h86;
	15'h130a: q<=8'h37;
	15'h130b: q<=8'ha9;
	15'h130c: q<=8'hff;
	15'h130d: q<=8'h9d;
	15'h130e: q<=8'hf2;
	15'h130f: q<=8'h02;
	15'h1310: q<=8'h98;
	15'h1311: q<=8'h38;
	15'h1312: q<=8'he9;
	15'h1313: q<=8'h04;
	15'h1314: q<=8'ha8;
	15'h1315: q<=8'hb9;
	15'h1316: q<=8'hb9;
	15'h1317: q<=8'h02;
	15'h1318: q<=8'h85;
	15'h1319: q<=8'h2d;
	15'h131a: q<=8'had;
	15'h131b: q<=8'hda;
	15'h131c: q<=8'h60;
	15'h131d: q<=8'h29;
	15'h131e: q<=8'h07;
	15'h131f: q<=8'hc9;
	15'h1320: q<=8'h03;
	15'h1321: q<=8'h90;
	15'h1322: q<=8'h02;
	15'h1323: q<=8'ha9;
	15'h1324: q<=8'h00;
	15'h1325: q<=8'h48;
	15'h1326: q<=8'h18;
	15'h1327: q<=8'h69;
	15'h1328: q<=8'h02;
	15'h1329: q<=8'h20;
	15'h132a: q<=8'hca;
	15'h132b: q<=8'ha3;
	15'h132c: q<=8'h20;
	15'h132d: q<=8'h6f;
	15'h132e: q<=8'ha0;
	15'h132f: q<=8'h68;
	15'h1330: q<=8'h18;
	15'h1331: q<=8'h69;
	15'h1332: q<=8'h05;
	15'h1333: q<=8'haa;
	15'h1334: q<=8'h20;
	15'h1335: q<=8'h6c;
	15'h1336: q<=8'hca;
	15'h1337: q<=8'ha6;
	15'h1338: q<=8'h37;
	15'h1339: q<=8'h60;
	15'h133a: q<=8'ha9;
	15'h133b: q<=8'h05;
	15'h133c: q<=8'h20;
	15'h133d: q<=8'h52;
	15'h133e: q<=8'ha3;
	15'h133f: q<=8'hce;
	15'h1340: q<=8'h01;
	15'h1341: q<=8'h02;
	15'h1342: q<=8'h60;
	15'h1343: q<=8'ha9;
	15'h1344: q<=8'h09;
	15'h1345: q<=8'hd0;
	15'h1346: q<=8'h06;
	15'h1347: q<=8'ha9;
	15'h1348: q<=8'h07;
	15'h1349: q<=8'hd0;
	15'h134a: q<=8'h02;
	15'h134b: q<=8'ha9;
	15'h134c: q<=8'hff;
	15'h134d: q<=8'h8d;
	15'h134e: q<=8'h3b;
	15'h134f: q<=8'h01;
	15'h1350: q<=8'ha9;
	15'h1351: q<=8'h01;
	15'h1352: q<=8'h85;
	15'h1353: q<=8'h2c;
	15'h1354: q<=8'had;
	15'h1355: q<=8'h02;
	15'h1356: q<=8'h02;
	15'h1357: q<=8'h85;
	15'h1358: q<=8'h29;
	15'h1359: q<=8'had;
	15'h135a: q<=8'h00;
	15'h135b: q<=8'h02;
	15'h135c: q<=8'h85;
	15'h135d: q<=8'h2d;
	15'h135e: q<=8'h20;
	15'h135f: q<=8'hb0;
	15'h1360: q<=8'hcc;
	15'h1361: q<=8'h20;
	15'h1362: q<=8'hd6;
	15'h1363: q<=8'ha3;
	15'h1364: q<=8'ha9;
	15'h1365: q<=8'h81;
	15'h1366: q<=8'h8d;
	15'h1367: q<=8'h01;
	15'h1368: q<=8'h02;
	15'h1369: q<=8'ha9;
	15'h136a: q<=8'h01;
	15'h136b: q<=8'h8d;
	15'h136c: q<=8'h3c;
	15'h136d: q<=8'h01;
	15'h136e: q<=8'h60;
	15'h136f: q<=8'h20;
	15'h1370: q<=8'hc1;
	15'h1371: q<=8'hcc;
	15'h1372: q<=8'hb9;
	15'h1373: q<=8'hdb;
	15'h1374: q<=8'h02;
	15'h1375: q<=8'h85;
	15'h1376: q<=8'h29;
	15'h1377: q<=8'hb9;
	15'h1378: q<=8'hb5;
	15'h1379: q<=8'h02;
	15'h137a: q<=8'h85;
	15'h137b: q<=8'h2d;
	15'h137c: q<=8'ha9;
	15'h137d: q<=8'h00;
	15'h137e: q<=8'h20;
	15'h137f: q<=8'hd4;
	15'h1380: q<=8'ha3;
	15'h1381: q<=8'ha9;
	15'h1382: q<=8'h00;
	15'h1383: q<=8'h99;
	15'h1384: q<=8'hdb;
	15'h1385: q<=8'h02;
	15'h1386: q<=8'hc6;
	15'h1387: q<=8'ha6;
	15'h1388: q<=8'ha9;
	15'h1389: q<=8'hff;
	15'h138a: q<=8'h9d;
	15'h138b: q<=8'hf2;
	15'h138c: q<=8'h02;
	15'h138d: q<=8'h60;
	15'h138e: q<=8'ha9;
	15'h138f: q<=8'hff;
	15'h1390: q<=8'h9d;
	15'h1391: q<=8'hf2;
	15'h1392: q<=8'h02;
	15'h1393: q<=8'h98;
	15'h1394: q<=8'h38;
	15'h1395: q<=8'he9;
	15'h1396: q<=8'h04;
	15'h1397: q<=8'ha8;
	15'h1398: q<=8'hb9;
	15'h1399: q<=8'h83;
	15'h139a: q<=8'h02;
	15'h139b: q<=8'h29;
	15'h139c: q<=8'hc0;
	15'h139d: q<=8'hc9;
	15'h139e: q<=8'hc0;
	15'h139f: q<=8'hf0;
	15'h13a0: q<=8'h06;
	15'h13a1: q<=8'hb9;
	15'h13a2: q<=8'hb9;
	15'h13a3: q<=8'h02;
	15'h13a4: q<=8'hb8;
	15'h13a5: q<=8'h50;
	15'h13a6: q<=8'h08;
	15'h13a7: q<=8'hb9;
	15'h13a8: q<=8'hb9;
	15'h13a9: q<=8'h02;
	15'h13aa: q<=8'h38;
	15'h13ab: q<=8'he9;
	15'h13ac: q<=8'h01;
	15'h13ad: q<=8'h29;
	15'h13ae: q<=8'h0f;
	15'h13af: q<=8'h85;
	15'h13b0: q<=8'h2d;
	15'h13b1: q<=8'ha9;
	15'h13b2: q<=8'h00;
	15'h13b3: q<=8'h20;
	15'h13b4: q<=8'hca;
	15'h13b5: q<=8'ha3;
	15'h13b6: q<=8'h20;
	15'h13b7: q<=8'h6f;
	15'h13b8: q<=8'ha0;
	15'h13b9: q<=8'hb9;
	15'h13ba: q<=8'h83;
	15'h13bb: q<=8'h02;
	15'h13bc: q<=8'h29;
	15'h13bd: q<=8'h07;
	15'h13be: q<=8'ha8;
	15'h13bf: q<=8'hbe;
	15'h13c0: q<=8'hc5;
	15'h13c1: q<=8'ha3;
	15'h13c2: q<=8'h4c;
	15'h13c3: q<=8'h6c;
	15'h13c4: q<=8'hca;
	15'h13c5: q<=8'h01;
	15'h13c6: q<=8'h02;
	15'h13c7: q<=8'h03;
	15'h13c8: q<=8'h04;
	15'h13c9: q<=8'h01;
	15'h13ca: q<=8'h48;
	15'h13cb: q<=8'h20;
	15'h13cc: q<=8'hc1;
	15'h13cd: q<=8'hcc;
	15'h13ce: q<=8'hb9;
	15'h13cf: q<=8'hdf;
	15'h13d0: q<=8'h02;
	15'h13d1: q<=8'h85;
	15'h13d2: q<=8'h29;
	15'h13d3: q<=8'h68;
	15'h13d4: q<=8'h85;
	15'h13d5: q<=8'h2c;
	15'h13d6: q<=8'h86;
	15'h13d7: q<=8'h35;
	15'h13d8: q<=8'h84;
	15'h13d9: q<=8'h36;
	15'h13da: q<=8'ha9;
	15'h13db: q<=8'h00;
	15'h13dc: q<=8'h85;
	15'h13dd: q<=8'h2a;
	15'h13de: q<=8'h85;
	15'h13df: q<=8'h2b;
	15'h13e0: q<=8'ha2;
	15'h13e1: q<=8'h07;
	15'h13e2: q<=8'hbd;
	15'h13e3: q<=8'h0a;
	15'h13e4: q<=8'h03;
	15'h13e5: q<=8'hf0;
	15'h13e6: q<=8'h13;
	15'h13e7: q<=8'hbd;
	15'h13e8: q<=8'h12;
	15'h13e9: q<=8'h03;
	15'h13ea: q<=8'hc5;
	15'h13eb: q<=8'h2a;
	15'h13ec: q<=8'h90;
	15'h13ed: q<=8'h04;
	15'h13ee: q<=8'h85;
	15'h13ef: q<=8'h2a;
	15'h13f0: q<=8'h86;
	15'h13f1: q<=8'h2b;
	15'h13f2: q<=8'hca;
	15'h13f3: q<=8'h10;
	15'h13f4: q<=8'hed;
	15'h13f5: q<=8'hce;
	15'h13f6: q<=8'h16;
	15'h13f7: q<=8'h01;
	15'h13f8: q<=8'ha6;
	15'h13f9: q<=8'h2b;
	15'h13fa: q<=8'ha9;
	15'h13fb: q<=8'h00;
	15'h13fc: q<=8'h9d;
	15'h13fd: q<=8'h12;
	15'h13fe: q<=8'h03;
	15'h13ff: q<=8'ha5;
	15'h1400: q<=8'h2c;
	15'h1401: q<=8'h9d;
	15'h1402: q<=8'h02;
	15'h1403: q<=8'h03;
	15'h1404: q<=8'ha5;
	15'h1405: q<=8'h29;
	15'h1406: q<=8'h9d;
	15'h1407: q<=8'h0a;
	15'h1408: q<=8'h03;
	15'h1409: q<=8'ha5;
	15'h140a: q<=8'h2d;
	15'h140b: q<=8'h9d;
	15'h140c: q<=8'hfa;
	15'h140d: q<=8'h02;
	15'h140e: q<=8'hee;
	15'h140f: q<=8'h16;
	15'h1410: q<=8'h01;
	15'h1411: q<=8'ha6;
	15'h1412: q<=8'h35;
	15'h1413: q<=8'ha4;
	15'h1414: q<=8'h36;
	15'h1415: q<=8'h60;
	15'h1416: q<=8'had;
	15'h1417: q<=8'h16;
	15'h1418: q<=8'h01;
	15'h1419: q<=8'hf0;
	15'h141a: q<=8'h2c;
	15'h141b: q<=8'ha9;
	15'h141c: q<=8'h00;
	15'h141d: q<=8'h8d;
	15'h141e: q<=8'h16;
	15'h141f: q<=8'h01;
	15'h1420: q<=8'ha2;
	15'h1421: q<=8'h07;
	15'h1422: q<=8'hbd;
	15'h1423: q<=8'h0a;
	15'h1424: q<=8'h03;
	15'h1425: q<=8'hf0;
	15'h1426: q<=8'h1d;
	15'h1427: q<=8'hbd;
	15'h1428: q<=8'h12;
	15'h1429: q<=8'h03;
	15'h142a: q<=8'hbc;
	15'h142b: q<=8'h02;
	15'h142c: q<=8'h03;
	15'h142d: q<=8'h18;
	15'h142e: q<=8'h79;
	15'h142f: q<=8'h4e;
	15'h1430: q<=8'ha4;
	15'h1431: q<=8'h9d;
	15'h1432: q<=8'h12;
	15'h1433: q<=8'h03;
	15'h1434: q<=8'hd9;
	15'h1435: q<=8'h48;
	15'h1436: q<=8'ha4;
	15'h1437: q<=8'h90;
	15'h1438: q<=8'h08;
	15'h1439: q<=8'ha9;
	15'h143a: q<=8'h00;
	15'h143b: q<=8'h9d;
	15'h143c: q<=8'h0a;
	15'h143d: q<=8'h03;
	15'h143e: q<=8'hb8;
	15'h143f: q<=8'h50;
	15'h1440: q<=8'h03;
	15'h1441: q<=8'hee;
	15'h1442: q<=8'h16;
	15'h1443: q<=8'h01;
	15'h1444: q<=8'hca;
	15'h1445: q<=8'h10;
	15'h1446: q<=8'hdb;
	15'h1447: q<=8'h60;
	15'h1448: q<=8'h10;
	15'h1449: q<=8'h15;
	15'h144a: q<=8'h20;
	15'h144b: q<=8'h20;
	15'h144c: q<=8'h20;
	15'h144d: q<=8'h10;
	15'h144e: q<=8'h03;
	15'h144f: q<=8'h01;
	15'h1450: q<=8'h03;
	15'h1451: q<=8'h03;
	15'h1452: q<=8'h03;
	15'h1453: q<=8'h03;
	15'h1454: q<=8'ha2;
	15'h1455: q<=8'h07;
	15'h1456: q<=8'hbd;
	15'h1457: q<=8'hd3;
	15'h1458: q<=8'h02;
	15'h1459: q<=8'hf0;
	15'h145a: q<=8'h03;
	15'h145b: q<=8'h20;
	15'h145c: q<=8'h63;
	15'h145d: q<=8'ha4;
	15'h145e: q<=8'hca;
	15'h145f: q<=8'h10;
	15'h1460: q<=8'hf5;
	15'h1461: q<=8'h60;
	15'h1462: q<=8'hab;
	15'h1463: q<=8'h85;
	15'h1464: q<=8'h2e;
	15'h1465: q<=8'ha0;
	15'h1466: q<=8'h0a;
	15'h1467: q<=8'hb9;
	15'h1468: q<=8'hdb;
	15'h1469: q<=8'h02;
	15'h146a: q<=8'hf0;
	15'h146b: q<=8'h7f;
	15'h146c: q<=8'hc5;
	15'h146d: q<=8'h2e;
	15'h146e: q<=8'h90;
	15'h146f: q<=8'h05;
	15'h1470: q<=8'he5;
	15'h1471: q<=8'h2e;
	15'h1472: q<=8'hb8;
	15'h1473: q<=8'h50;
	15'h1474: q<=8'h06;
	15'h1475: q<=8'ha5;
	15'h1476: q<=8'h2e;
	15'h1477: q<=8'h38;
	15'h1478: q<=8'hf9;
	15'h1479: q<=8'hdb;
	15'h147a: q<=8'h02;
	15'h147b: q<=8'hc0;
	15'h147c: q<=8'h04;
	15'h147d: q<=8'hb0;
	15'h147e: q<=8'h12;
	15'h147f: q<=8'hc5;
	15'h1480: q<=8'ha7;
	15'h1481: q<=8'hb0;
	15'h1482: q<=8'h0b;
	15'h1483: q<=8'hb9;
	15'h1484: q<=8'hb5;
	15'h1485: q<=8'h02;
	15'h1486: q<=8'h5d;
	15'h1487: q<=8'had;
	15'h1488: q<=8'h02;
	15'h1489: q<=8'hd0;
	15'h148a: q<=8'h03;
	15'h148b: q<=8'h20;
	15'h148c: q<=8'h6f;
	15'h148d: q<=8'ha3;
	15'h148e: q<=8'hb8;
	15'h148f: q<=8'h50;
	15'h1490: q<=8'h5a;
	15'h1491: q<=8'h48;
	15'h1492: q<=8'h84;
	15'h1493: q<=8'h38;
	15'h1494: q<=8'hb9;
	15'h1495: q<=8'h7f;
	15'h1496: q<=8'h02;
	15'h1497: q<=8'h29;
	15'h1498: q<=8'h07;
	15'h1499: q<=8'ha8;
	15'h149a: q<=8'h68;
	15'h149b: q<=8'hd9;
	15'h149c: q<=8'h51;
	15'h149d: q<=8'h01;
	15'h149e: q<=8'hb0;
	15'h149f: q<=8'h49;
	15'h14a0: q<=8'hc0;
	15'h14a1: q<=8'h04;
	15'h14a2: q<=8'hd0;
	15'h14a3: q<=8'h1d;
	15'h14a4: q<=8'ha4;
	15'h14a5: q<=8'h38;
	15'h14a6: q<=8'hb9;
	15'h14a7: q<=8'hdb;
	15'h14a8: q<=8'h02;
	15'h14a9: q<=8'hcd;
	15'h14aa: q<=8'h02;
	15'h14ab: q<=8'h02;
	15'h14ac: q<=8'hf0;
	15'h14ad: q<=8'h10;
	15'h14ae: q<=8'hbd;
	15'h14af: q<=8'had;
	15'h14b0: q<=8'h02;
	15'h14b1: q<=8'hd9;
	15'h14b2: q<=8'hb5;
	15'h14b3: q<=8'h02;
	15'h14b4: q<=8'hd0;
	15'h14b5: q<=8'h08;
	15'h14b6: q<=8'hb9;
	15'h14b7: q<=8'hc8;
	15'h14b8: q<=8'h02;
	15'h14b9: q<=8'h10;
	15'h14ba: q<=8'h03;
	15'h14bb: q<=8'h20;
	15'h14bc: q<=8'h09;
	15'h14bd: q<=8'ha3;
	15'h14be: q<=8'hb8;
	15'h14bf: q<=8'h50;
	15'h14c0: q<=8'h28;
	15'h14c1: q<=8'ha4;
	15'h14c2: q<=8'h38;
	15'h14c3: q<=8'hb9;
	15'h14c4: q<=8'hc8;
	15'h14c5: q<=8'h02;
	15'h14c6: q<=8'h10;
	15'h14c7: q<=8'h0a;
	15'h14c8: q<=8'hb9;
	15'h14c9: q<=8'hb5;
	15'h14ca: q<=8'h02;
	15'h14cb: q<=8'hdd;
	15'h14cc: q<=8'hc0;
	15'h14cd: q<=8'h02;
	15'h14ce: q<=8'hf0;
	15'h14cf: q<=8'h12;
	15'h14d0: q<=8'hd0;
	15'h14d1: q<=8'h08;
	15'h14d2: q<=8'hb9;
	15'h14d3: q<=8'hdb;
	15'h14d4: q<=8'h02;
	15'h14d5: q<=8'hcd;
	15'h14d6: q<=8'h02;
	15'h14d7: q<=8'h02;
	15'h14d8: q<=8'hf0;
	15'h14d9: q<=8'h0f;
	15'h14da: q<=8'hb9;
	15'h14db: q<=8'hb5;
	15'h14dc: q<=8'h02;
	15'h14dd: q<=8'hdd;
	15'h14de: q<=8'had;
	15'h14df: q<=8'h02;
	15'h14e0: q<=8'hd0;
	15'h14e1: q<=8'h07;
	15'h14e2: q<=8'h86;
	15'h14e3: q<=8'h37;
	15'h14e4: q<=8'h20;
	15'h14e5: q<=8'h8e;
	15'h14e6: q<=8'ha3;
	15'h14e7: q<=8'ha6;
	15'h14e8: q<=8'h37;
	15'h14e9: q<=8'ha4;
	15'h14ea: q<=8'h38;
	15'h14eb: q<=8'h88;
	15'h14ec: q<=8'h30;
	15'h14ed: q<=8'h03;
	15'h14ee: q<=8'h4c;
	15'h14ef: q<=8'h67;
	15'h14f0: q<=8'ha4;
	15'h14f1: q<=8'hbd;
	15'h14f2: q<=8'hf2;
	15'h14f3: q<=8'h02;
	15'h14f4: q<=8'hc9;
	15'h14f5: q<=8'hff;
	15'h14f6: q<=8'hd0;
	15'h14f7: q<=8'h0b;
	15'h14f8: q<=8'ha9;
	15'h14f9: q<=8'h00;
	15'h14fa: q<=8'h9d;
	15'h14fb: q<=8'hd3;
	15'h14fc: q<=8'h02;
	15'h14fd: q<=8'hce;
	15'h14fe: q<=8'h35;
	15'h14ff: q<=8'h01;
	15'h1500: q<=8'h9d;
	15'h1501: q<=8'hf2;
	15'h1502: q<=8'h02;
	15'h1503: q<=8'h60;
	15'h1504: q<=8'had;
	15'h1505: q<=8'h01;
	15'h1506: q<=8'h02;
	15'h1507: q<=8'h10;
	15'h1508: q<=8'h78;
	15'h1509: q<=8'had;
	15'h150a: q<=8'h35;
	15'h150b: q<=8'h01;
	15'h150c: q<=8'h05;
	15'h150d: q<=8'ha6;
	15'h150e: q<=8'h0d;
	15'h150f: q<=8'h16;
	15'h1510: q<=8'h01;
	15'h1511: q<=8'hd0;
	15'h1512: q<=8'h6b;
	15'h1513: q<=8'hae;
	15'h1514: q<=8'h1c;
	15'h1515: q<=8'h01;
	15'h1516: q<=8'hbd;
	15'h1517: q<=8'hdf;
	15'h1518: q<=8'h02;
	15'h1519: q<=8'hf0;
	15'h151a: q<=8'h0e;
	15'h151b: q<=8'h18;
	15'h151c: q<=8'h69;
	15'h151d: q<=8'h0f;
	15'h151e: q<=8'hb0;
	15'h151f: q<=8'h02;
	15'h1520: q<=8'hc9;
	15'h1521: q<=8'hf0;
	15'h1522: q<=8'h90;
	15'h1523: q<=8'h02;
	15'h1524: q<=8'ha9;
	15'h1525: q<=8'h00;
	15'h1526: q<=8'h9d;
	15'h1527: q<=8'hdf;
	15'h1528: q<=8'h02;
	15'h1529: q<=8'hca;
	15'h152a: q<=8'h10;
	15'h152b: q<=8'hea;
	15'h152c: q<=8'ha6;
	15'h152d: q<=8'h3d;
	15'h152e: q<=8'hb5;
	15'h152f: q<=8'h48;
	15'h1530: q<=8'hc9;
	15'h1531: q<=8'h01;
	15'h1532: q<=8'hd0;
	15'h1533: q<=8'h20;
	15'h1534: q<=8'ha9;
	15'h1535: q<=8'h00;
	15'h1536: q<=8'h8d;
	15'h1537: q<=8'h0f;
	15'h1538: q<=8'h01;
	15'h1539: q<=8'ha9;
	15'h153a: q<=8'h01;
	15'h153b: q<=8'h8d;
	15'h153c: q<=8'h14;
	15'h153d: q<=8'h01;
	15'h153e: q<=8'ha5;
	15'h153f: q<=8'h5f;
	15'h1540: q<=8'h38;
	15'h1541: q<=8'he9;
	15'h1542: q<=8'h20;
	15'h1543: q<=8'h85;
	15'h1544: q<=8'h5f;
	15'h1545: q<=8'ha5;
	15'h1546: q<=8'h5b;
	15'h1547: q<=8'he9;
	15'h1548: q<=8'h00;
	15'h1549: q<=8'h85;
	15'h154a: q<=8'h5b;
	15'h154b: q<=8'hc9;
	15'h154c: q<=8'hfa;
	15'h154d: q<=8'h18;
	15'h154e: q<=8'hd0;
	15'h154f: q<=8'h01;
	15'h1550: q<=8'h38;
	15'h1551: q<=8'hb8;
	15'h1552: q<=8'h50;
	15'h1553: q<=8'h0d;
	15'h1554: q<=8'had;
	15'h1555: q<=8'h02;
	15'h1556: q<=8'h02;
	15'h1557: q<=8'h18;
	15'h1558: q<=8'h69;
	15'h1559: q<=8'h0f;
	15'h155a: q<=8'h8d;
	15'h155b: q<=8'h02;
	15'h155c: q<=8'h02;
	15'h155d: q<=8'hb0;
	15'h155e: q<=8'h02;
	15'h155f: q<=8'hc9;
	15'h1560: q<=8'hf0;
	15'h1561: q<=8'h90;
	15'h1562: q<=8'h1b;
	15'h1563: q<=8'ha9;
	15'h1564: q<=8'h06;
	15'h1565: q<=8'h85;
	15'h1566: q<=8'h00;
	15'h1567: q<=8'h20;
	15'h1568: q<=8'h8f;
	15'h1569: q<=8'h92;
	15'h156a: q<=8'had;
	15'h156b: q<=8'h08;
	15'h156c: q<=8'h01;
	15'h156d: q<=8'h18;
	15'h156e: q<=8'h6d;
	15'h156f: q<=8'h09;
	15'h1570: q<=8'h01;
	15'h1571: q<=8'h18;
	15'h1572: q<=8'h6d;
	15'h1573: q<=8'hab;
	15'h1574: q<=8'h03;
	15'h1575: q<=8'hc9;
	15'h1576: q<=8'h3f;
	15'h1577: q<=8'h90;
	15'h1578: q<=8'h02;
	15'h1579: q<=8'ha9;
	15'h157a: q<=8'h3f;
	15'h157b: q<=8'h8d;
	15'h157c: q<=8'hab;
	15'h157d: q<=8'h03;
	15'h157e: q<=8'hb8;
	15'h157f: q<=8'h50;
	15'h1580: q<=8'h49;
	15'h1581: q<=8'had;
	15'h1582: q<=8'h55;
	15'h1583: q<=8'h04;
	15'h1584: q<=8'h0d;
	15'h1585: q<=8'h1b;
	15'h1586: q<=8'h01;
	15'h1587: q<=8'hf0;
	15'h1588: q<=8'h0a;
	15'h1589: q<=8'ha9;
	15'h158a: q<=8'h17;
	15'h158b: q<=8'hc5;
	15'h158c: q<=8'h42;
	15'h158d: q<=8'hb0;
	15'h158e: q<=8'h04;
	15'h158f: q<=8'ha6;
	15'h1590: q<=8'h40;
	15'h1591: q<=8'hf6;
	15'h1592: q<=8'h00;
	15'h1593: q<=8'had;
	15'h1594: q<=8'h06;
	15'h1595: q<=8'h01;
	15'h1596: q<=8'hd0;
	15'h1597: q<=8'h32;
	15'h1598: q<=8'had;
	15'h1599: q<=8'hab;
	15'h159a: q<=8'h03;
	15'h159b: q<=8'h0d;
	15'h159c: q<=8'h16;
	15'h159d: q<=8'h01;
	15'h159e: q<=8'hd0;
	15'h159f: q<=8'h15;
	15'h15a0: q<=8'hac;
	15'h15a1: q<=8'h1c;
	15'h15a2: q<=8'h01;
	15'h15a3: q<=8'hb9;
	15'h15a4: q<=8'hdf;
	15'h15a5: q<=8'h02;
	15'h15a6: q<=8'hf0;
	15'h15a7: q<=8'h04;
	15'h15a8: q<=8'hc9;
	15'h15a9: q<=8'h11;
	15'h15aa: q<=8'hb0;
	15'h15ab: q<=8'h09;
	15'h15ac: q<=8'h88;
	15'h15ad: q<=8'h10;
	15'h15ae: q<=8'hf4;
	15'h15af: q<=8'h20;
	15'h15b0: q<=8'hcb;
	15'h15b1: q<=8'ha5;
	15'h15b2: q<=8'h20;
	15'h15b3: q<=8'h8f;
	15'h15b4: q<=8'h92;
	15'h15b5: q<=8'ha5;
	15'h15b6: q<=8'h4d;
	15'h15b7: q<=8'h29;
	15'h15b8: q<=8'h60;
	15'h15b9: q<=8'hf0;
	15'h15ba: q<=8'h0f;
	15'h15bb: q<=8'h24;
	15'h15bc: q<=8'h05;
	15'h15bd: q<=8'h10;
	15'h15be: q<=8'h0b;
	15'h15bf: q<=8'ha5;
	15'h15c0: q<=8'h09;
	15'h15c1: q<=8'h29;
	15'h15c2: q<=8'h43;
	15'h15c3: q<=8'hc9;
	15'h15c4: q<=8'h40;
	15'h15c5: q<=8'hd0;
	15'h15c6: q<=8'h03;
	15'h15c7: q<=8'h20;
	15'h15c8: q<=8'hcb;
	15'h15c9: q<=8'ha5;
	15'h15ca: q<=8'h60;
	15'h15cb: q<=8'ha9;
	15'h15cc: q<=8'h20;
	15'h15cd: q<=8'h85;
	15'h15ce: q<=8'h00;
	15'h15cf: q<=8'had;
	15'h15d0: q<=8'h06;
	15'h15d1: q<=8'h01;
	15'h15d2: q<=8'h09;
	15'h15d3: q<=8'h80;
	15'h15d4: q<=8'h8d;
	15'h15d5: q<=8'h06;
	15'h15d6: q<=8'h01;
	15'h15d7: q<=8'ha9;
	15'h15d8: q<=8'h00;
	15'h15d9: q<=8'h8d;
	15'h15da: q<=8'h04;
	15'h15db: q<=8'h01;
	15'h15dc: q<=8'h8d;
	15'h15dd: q<=8'h07;
	15'h15de: q<=8'h01;
	15'h15df: q<=8'h85;
	15'h15e0: q<=8'h5c;
	15'h15e1: q<=8'h8d;
	15'h15e2: q<=8'h23;
	15'h15e3: q<=8'h01;
	15'h15e4: q<=8'ha9;
	15'h15e5: q<=8'h02;
	15'h15e6: q<=8'h8d;
	15'h15e7: q<=8'h05;
	15'h15e8: q<=8'h01;
	15'h15e9: q<=8'ha2;
	15'h15ea: q<=8'h0f;
	15'h15eb: q<=8'hbd;
	15'h15ec: q<=8'hac;
	15'h15ed: q<=8'h03;
	15'h15ee: q<=8'hf0;
	15'h15ef: q<=8'h03;
	15'h15f0: q<=8'hee;
	15'h15f1: q<=8'h23;
	15'h15f2: q<=8'h01;
	15'h15f3: q<=8'hca;
	15'h15f4: q<=8'h10;
	15'h15f5: q<=8'hf5;
	15'h15f6: q<=8'had;
	15'h15f7: q<=8'h23;
	15'h15f8: q<=8'h01;
	15'h15f9: q<=8'hf0;
	15'h15fa: q<=8'h17;
	15'h15fb: q<=8'ha5;
	15'h15fc: q<=8'h9f;
	15'h15fd: q<=8'hc9;
	15'h15fe: q<=8'h07;
	15'h15ff: q<=8'hb0;
	15'h1600: q<=8'h11;
	15'h1601: q<=8'ha9;
	15'h1602: q<=8'h1e;
	15'h1603: q<=8'h85;
	15'h1604: q<=8'h04;
	15'h1605: q<=8'ha9;
	15'h1606: q<=8'h0a;
	15'h1607: q<=8'h85;
	15'h1608: q<=8'h00;
	15'h1609: q<=8'ha9;
	15'h160a: q<=8'h20;
	15'h160b: q<=8'h85;
	15'h160c: q<=8'h02;
	15'h160d: q<=8'ha9;
	15'h160e: q<=8'h80;
	15'h160f: q<=8'h8d;
	15'h1610: q<=8'h23;
	15'h1611: q<=8'h01;
	15'h1612: q<=8'ha9;
	15'h1613: q<=8'hff;
	15'h1614: q<=8'h8d;
	15'h1615: q<=8'h25;
	15'h1616: q<=8'h01;
	15'h1617: q<=8'h60;
	15'h1618: q<=8'had;
	15'h1619: q<=8'h0e;
	15'h161a: q<=8'h01;
	15'h161b: q<=8'h8d;
	15'h161c: q<=8'h0d;
	15'h161d: q<=8'h01;
	15'h161e: q<=8'ha2;
	15'h161f: q<=8'h0f;
	15'h1620: q<=8'h86;
	15'h1621: q<=8'h37;
	15'h1622: q<=8'ha6;
	15'h1623: q<=8'h37;
	15'h1624: q<=8'hbd;
	15'h1625: q<=8'h83;
	15'h1626: q<=8'h02;
	15'h1627: q<=8'hd0;
	15'h1628: q<=8'h0b;
	15'h1629: q<=8'had;
	15'h162a: q<=8'h0e;
	15'h162b: q<=8'h01;
	15'h162c: q<=8'hf0;
	15'h162d: q<=8'h03;
	15'h162e: q<=8'h20;
	15'h162f: q<=8'h5b;
	15'h1630: q<=8'ha6;
	15'h1631: q<=8'hb8;
	15'h1632: q<=8'h50;
	15'h1633: q<=8'h0b;
	15'h1634: q<=8'h20;
	15'h1635: q<=8'ha9;
	15'h1636: q<=8'ha6;
	15'h1637: q<=8'h20;
	15'h1638: q<=8'h21;
	15'h1639: q<=8'ha7;
	15'h163a: q<=8'ha9;
	15'h163b: q<=8'hff;
	15'h163c: q<=8'h8d;
	15'h163d: q<=8'h0d;
	15'h163e: q<=8'h01;
	15'h163f: q<=8'hc6;
	15'h1640: q<=8'h37;
	15'h1641: q<=8'h10;
	15'h1642: q<=8'hdf;
	15'h1643: q<=8'ha5;
	15'h1644: q<=8'h03;
	15'h1645: q<=8'h29;
	15'h1646: q<=8'h01;
	15'h1647: q<=8'hd0;
	15'h1648: q<=8'h08;
	15'h1649: q<=8'had;
	15'h164a: q<=8'h0e;
	15'h164b: q<=8'h01;
	15'h164c: q<=8'hf0;
	15'h164d: q<=8'h03;
	15'h164e: q<=8'hce;
	15'h164f: q<=8'h0e;
	15'h1650: q<=8'h01;
	15'h1651: q<=8'had;
	15'h1652: q<=8'h0d;
	15'h1653: q<=8'h01;
	15'h1654: q<=8'hd0;
	15'h1655: q<=8'h04;
	15'h1656: q<=8'ha9;
	15'h1657: q<=8'h12;
	15'h1658: q<=8'h85;
	15'h1659: q<=8'h00;
	15'h165a: q<=8'h60;
	15'h165b: q<=8'ha5;
	15'h165c: q<=8'h03;
	15'h165d: q<=8'h29;
	15'h165e: q<=8'h00;
	15'h165f: q<=8'hd0;
	15'h1660: q<=8'h39;
	15'h1661: q<=8'ha9;
	15'h1662: q<=8'h80;
	15'h1663: q<=8'h9d;
	15'h1664: q<=8'h63;
	15'h1665: q<=8'h02;
	15'h1666: q<=8'h9d;
	15'h1667: q<=8'h83;
	15'h1668: q<=8'h02;
	15'h1669: q<=8'h9d;
	15'h166a: q<=8'ha3;
	15'h166b: q<=8'h02;
	15'h166c: q<=8'had;
	15'h166d: q<=8'hda;
	15'h166e: q<=8'h60;
	15'h166f: q<=8'h9d;
	15'h1670: q<=8'hc3;
	15'h1671: q<=8'h02;
	15'h1672: q<=8'h20;
	15'h1673: q<=8'h9b;
	15'h1674: q<=8'ha6;
	15'h1675: q<=8'h9d;
	15'h1676: q<=8'h23;
	15'h1677: q<=8'h03;
	15'h1678: q<=8'had;
	15'h1679: q<=8'hca;
	15'h167a: q<=8'h60;
	15'h167b: q<=8'h9d;
	15'h167c: q<=8'he3;
	15'h167d: q<=8'h02;
	15'h167e: q<=8'h20;
	15'h167f: q<=8'h9b;
	15'h1680: q<=8'ha6;
	15'h1681: q<=8'h30;
	15'h1682: q<=8'h05;
	15'h1683: q<=8'h49;
	15'h1684: q<=8'hff;
	15'h1685: q<=8'h18;
	15'h1686: q<=8'h69;
	15'h1687: q<=8'h01;
	15'h1688: q<=8'h9d;
	15'h1689: q<=8'h43;
	15'h168a: q<=8'h03;
	15'h168b: q<=8'had;
	15'h168c: q<=8'hca;
	15'h168d: q<=8'h60;
	15'h168e: q<=8'h9d;
	15'h168f: q<=8'h03;
	15'h1690: q<=8'h03;
	15'h1691: q<=8'h20;
	15'h1692: q<=8'h9b;
	15'h1693: q<=8'ha6;
	15'h1694: q<=8'h9d;
	15'h1695: q<=8'h63;
	15'h1696: q<=8'h03;
	15'h1697: q<=8'h20;
	15'h1698: q<=8'hc1;
	15'h1699: q<=8'hcc;
	15'h169a: q<=8'h60;
	15'h169b: q<=8'h4a;
	15'h169c: q<=8'had;
	15'h169d: q<=8'hda;
	15'h169e: q<=8'h60;
	15'h169f: q<=8'h29;
	15'h16a0: q<=8'h07;
	15'h16a1: q<=8'h90;
	15'h16a2: q<=8'h05;
	15'h16a3: q<=8'h49;
	15'h16a4: q<=8'hff;
	15'h16a5: q<=8'h18;
	15'h16a6: q<=8'h69;
	15'h16a7: q<=8'h01;
	15'h16a8: q<=8'h60;
	15'h16a9: q<=8'hbd;
	15'h16aa: q<=8'he3;
	15'h16ab: q<=8'h02;
	15'h16ac: q<=8'h18;
	15'h16ad: q<=8'h7d;
	15'h16ae: q<=8'h23;
	15'h16af: q<=8'h02;
	15'h16b0: q<=8'h9d;
	15'h16b1: q<=8'h23;
	15'h16b2: q<=8'h02;
	15'h16b3: q<=8'hbd;
	15'h16b4: q<=8'h43;
	15'h16b5: q<=8'h03;
	15'h16b6: q<=8'h30;
	15'h16b7: q<=8'h0c;
	15'h16b8: q<=8'h7d;
	15'h16b9: q<=8'h83;
	15'h16ba: q<=8'h02;
	15'h16bb: q<=8'hc9;
	15'h16bc: q<=8'hf0;
	15'h16bd: q<=8'h90;
	15'h16be: q<=8'h02;
	15'h16bf: q<=8'ha9;
	15'h16c0: q<=8'h00;
	15'h16c1: q<=8'hb8;
	15'h16c2: q<=8'h50;
	15'h16c3: q<=8'h09;
	15'h16c4: q<=8'h7d;
	15'h16c5: q<=8'h83;
	15'h16c6: q<=8'h02;
	15'h16c7: q<=8'hc9;
	15'h16c8: q<=8'h10;
	15'h16c9: q<=8'hb0;
	15'h16ca: q<=8'h02;
	15'h16cb: q<=8'ha9;
	15'h16cc: q<=8'h00;
	15'h16cd: q<=8'ha8;
	15'h16ce: q<=8'hbd;
	15'h16cf: q<=8'hc3;
	15'h16d0: q<=8'h02;
	15'h16d1: q<=8'h18;
	15'h16d2: q<=8'h7d;
	15'h16d3: q<=8'h03;
	15'h16d4: q<=8'h02;
	15'h16d5: q<=8'h9d;
	15'h16d6: q<=8'h03;
	15'h16d7: q<=8'h02;
	15'h16d8: q<=8'hbd;
	15'h16d9: q<=8'h23;
	15'h16da: q<=8'h03;
	15'h16db: q<=8'h30;
	15'h16dc: q<=8'h0c;
	15'h16dd: q<=8'h7d;
	15'h16de: q<=8'h63;
	15'h16df: q<=8'h02;
	15'h16e0: q<=8'hc9;
	15'h16e1: q<=8'hf0;
	15'h16e2: q<=8'h90;
	15'h16e3: q<=8'h02;
	15'h16e4: q<=8'ha0;
	15'h16e5: q<=8'h00;
	15'h16e6: q<=8'hb8;
	15'h16e7: q<=8'h50;
	15'h16e8: q<=8'h09;
	15'h16e9: q<=8'h7d;
	15'h16ea: q<=8'h63;
	15'h16eb: q<=8'h02;
	15'h16ec: q<=8'hc9;
	15'h16ed: q<=8'h10;
	15'h16ee: q<=8'hb0;
	15'h16ef: q<=8'h02;
	15'h16f0: q<=8'ha0;
	15'h16f1: q<=8'h00;
	15'h16f2: q<=8'h9d;
	15'h16f3: q<=8'h63;
	15'h16f4: q<=8'h02;
	15'h16f5: q<=8'hbd;
	15'h16f6: q<=8'h03;
	15'h16f7: q<=8'h03;
	15'h16f8: q<=8'h18;
	15'h16f9: q<=8'h7d;
	15'h16fa: q<=8'h43;
	15'h16fb: q<=8'h02;
	15'h16fc: q<=8'h9d;
	15'h16fd: q<=8'h43;
	15'h16fe: q<=8'h02;
	15'h16ff: q<=8'hbd;
	15'h1700: q<=8'h63;
	15'h1701: q<=8'h03;
	15'h1702: q<=8'h30;
	15'h1703: q<=8'h0c;
	15'h1704: q<=8'h7d;
	15'h1705: q<=8'ha3;
	15'h1706: q<=8'h02;
	15'h1707: q<=8'hc9;
	15'h1708: q<=8'hf0;
	15'h1709: q<=8'h90;
	15'h170a: q<=8'h02;
	15'h170b: q<=8'ha0;
	15'h170c: q<=8'h00;
	15'h170d: q<=8'hb8;
	15'h170e: q<=8'h50;
	15'h170f: q<=8'h09;
	15'h1710: q<=8'h7d;
	15'h1711: q<=8'ha3;
	15'h1712: q<=8'h02;
	15'h1713: q<=8'hc9;
	15'h1714: q<=8'h10;
	15'h1715: q<=8'hb0;
	15'h1716: q<=8'h02;
	15'h1717: q<=8'ha0;
	15'h1718: q<=8'h00;
	15'h1719: q<=8'h9d;
	15'h171a: q<=8'ha3;
	15'h171b: q<=8'h02;
	15'h171c: q<=8'h98;
	15'h171d: q<=8'h9d;
	15'h171e: q<=8'h83;
	15'h171f: q<=8'h02;
	15'h1720: q<=8'h60;
	15'h1721: q<=8'ha9;
	15'h1722: q<=8'hfd;
	15'h1723: q<=8'h85;
	15'h1724: q<=8'h29;
	15'h1725: q<=8'hbd;
	15'h1726: q<=8'hc3;
	15'h1727: q<=8'h02;
	15'h1728: q<=8'hbc;
	15'h1729: q<=8'h23;
	15'h172a: q<=8'h03;
	15'h172b: q<=8'h20;
	15'h172c: q<=8'h5d;
	15'h172d: q<=8'ha7;
	15'h172e: q<=8'h9d;
	15'h172f: q<=8'hc3;
	15'h1730: q<=8'h02;
	15'h1731: q<=8'h98;
	15'h1732: q<=8'h9d;
	15'h1733: q<=8'h23;
	15'h1734: q<=8'h03;
	15'h1735: q<=8'hbd;
	15'h1736: q<=8'he3;
	15'h1737: q<=8'h02;
	15'h1738: q<=8'hbc;
	15'h1739: q<=8'h43;
	15'h173a: q<=8'h03;
	15'h173b: q<=8'h20;
	15'h173c: q<=8'h5d;
	15'h173d: q<=8'ha7;
	15'h173e: q<=8'h9d;
	15'h173f: q<=8'he3;
	15'h1740: q<=8'h02;
	15'h1741: q<=8'h98;
	15'h1742: q<=8'h9d;
	15'h1743: q<=8'h43;
	15'h1744: q<=8'h03;
	15'h1745: q<=8'hbd;
	15'h1746: q<=8'h03;
	15'h1747: q<=8'h03;
	15'h1748: q<=8'hbc;
	15'h1749: q<=8'h63;
	15'h174a: q<=8'h03;
	15'h174b: q<=8'h20;
	15'h174c: q<=8'h5d;
	15'h174d: q<=8'ha7;
	15'h174e: q<=8'h9d;
	15'h174f: q<=8'h03;
	15'h1750: q<=8'h03;
	15'h1751: q<=8'h98;
	15'h1752: q<=8'h9d;
	15'h1753: q<=8'h63;
	15'h1754: q<=8'h03;
	15'h1755: q<=8'ha5;
	15'h1756: q<=8'h29;
	15'h1757: q<=8'hd0;
	15'h1758: q<=8'h03;
	15'h1759: q<=8'h9d;
	15'h175a: q<=8'h83;
	15'h175b: q<=8'h02;
	15'h175c: q<=8'h60;
	15'h175d: q<=8'h84;
	15'h175e: q<=8'h2b;
	15'h175f: q<=8'h24;
	15'h1760: q<=8'h2b;
	15'h1761: q<=8'h30;
	15'h1762: q<=8'h0f;
	15'h1763: q<=8'h38;
	15'h1764: q<=8'hed;
	15'h1765: q<=8'h88;
	15'h1766: q<=8'ha7;
	15'h1767: q<=8'h85;
	15'h1768: q<=8'h2a;
	15'h1769: q<=8'ha5;
	15'h176a: q<=8'h2b;
	15'h176b: q<=8'he9;
	15'h176c: q<=8'h00;
	15'h176d: q<=8'h90;
	15'h176e: q<=8'h0f;
	15'h176f: q<=8'hb8;
	15'h1770: q<=8'h50;
	15'h1771: q<=8'h12;
	15'h1772: q<=8'h18;
	15'h1773: q<=8'h6d;
	15'h1774: q<=8'h88;
	15'h1775: q<=8'ha7;
	15'h1776: q<=8'h85;
	15'h1777: q<=8'h2a;
	15'h1778: q<=8'ha5;
	15'h1779: q<=8'h2b;
	15'h177a: q<=8'h69;
	15'h177b: q<=8'h00;
	15'h177c: q<=8'h90;
	15'h177d: q<=8'h06;
	15'h177e: q<=8'he6;
	15'h177f: q<=8'h29;
	15'h1780: q<=8'ha9;
	15'h1781: q<=8'h00;
	15'h1782: q<=8'h85;
	15'h1783: q<=8'h2a;
	15'h1784: q<=8'ha8;
	15'h1785: q<=8'ha5;
	15'h1786: q<=8'h2a;
	15'h1787: q<=8'h60;
	15'h1788: q<=8'h20;
	15'h1789: q<=8'ha2;
	15'h178a: q<=8'h0f;
	15'h178b: q<=8'ha9;
	15'h178c: q<=8'h00;
	15'h178d: q<=8'h9d;
	15'h178e: q<=8'h83;
	15'h178f: q<=8'h02;
	15'h1790: q<=8'hca;
	15'h1791: q<=8'h10;
	15'h1792: q<=8'hf8;
	15'h1793: q<=8'ha9;
	15'h1794: q<=8'h20;
	15'h1795: q<=8'h8d;
	15'h1796: q<=8'h0e;
	15'h1797: q<=8'h01;
	15'h1798: q<=8'h8d;
	15'h1799: q<=8'h0d;
	15'h179a: q<=8'h01;
	15'h179b: q<=8'ha9;
	15'h179c: q<=8'h04;
	15'h179d: q<=8'h85;
	15'h179e: q<=8'h01;
	15'h179f: q<=8'ha9;
	15'h17a0: q<=8'h00;
	15'h17a1: q<=8'h85;
	15'h17a2: q<=8'h68;
	15'h17a3: q<=8'h85;
	15'h17a4: q<=8'h69;
	15'h17a5: q<=8'h60;
	15'h17a6: q<=8'h84;
	15'h17a7: q<=8'h2a;
	15'h17a8: q<=8'h38;
	15'h17a9: q<=8'he5;
	15'h17aa: q<=8'h2a;
	15'h17ab: q<=8'h85;
	15'h17ac: q<=8'h2a;
	15'h17ad: q<=8'h2c;
	15'h17ae: q<=8'h11;
	15'h17af: q<=8'h01;
	15'h17b0: q<=8'h30;
	15'h17b1: q<=8'h09;
	15'h17b2: q<=8'h29;
	15'h17b3: q<=8'h0f;
	15'h17b4: q<=8'h2c;
	15'h17b5: q<=8'hbc;
	15'h17b6: q<=8'ha7;
	15'h17b7: q<=8'hf0;
	15'h17b8: q<=8'h02;
	15'h17b9: q<=8'h09;
	15'h17ba: q<=8'hf8;
	15'h17bb: q<=8'h60;
	15'h17bc: q<=8'h08;
	15'h17bd: q<=8'ha2;
	15'h17be: q<=8'h07;
	15'h17bf: q<=8'ha9;
	15'h17c0: q<=8'h00;
	15'h17c1: q<=8'h9d;
	15'h17c2: q<=8'hfe;
	15'h17c3: q<=8'h03;
	15'h17c4: q<=8'hca;
	15'h17c5: q<=8'h10;
	15'h17c6: q<=8'hfa;
	15'h17c7: q<=8'ha9;
	15'h17c8: q<=8'hf0;
	15'h17c9: q<=8'h8d;
	15'h17ca: q<=8'h05;
	15'h17cb: q<=8'h04;
	15'h17cc: q<=8'ha9;
	15'h17cd: q<=8'hff;
	15'h17ce: q<=8'h8d;
	15'h17cf: q<=8'h15;
	15'h17d0: q<=8'h01;
	15'h17d1: q<=8'h60;
	15'h17d2: q<=8'had;
	15'h17d3: q<=8'h15;
	15'h17d4: q<=8'h01;
	15'h17d5: q<=8'hf0;
	15'h17d6: q<=8'h59;
	15'h17d7: q<=8'ha9;
	15'h17d8: q<=8'h00;
	15'h17d9: q<=8'h85;
	15'h17da: q<=8'h29;
	15'h17db: q<=8'ha2;
	15'h17dc: q<=8'h07;
	15'h17dd: q<=8'h86;
	15'h17de: q<=8'h37;
	15'h17df: q<=8'ha6;
	15'h17e0: q<=8'h37;
	15'h17e1: q<=8'hbd;
	15'h17e2: q<=8'hfe;
	15'h17e3: q<=8'h03;
	15'h17e4: q<=8'hf0;
	15'h17e5: q<=8'h18;
	15'h17e6: q<=8'h38;
	15'h17e7: q<=8'he9;
	15'h17e8: q<=8'h07;
	15'h17e9: q<=8'h90;
	15'h17ea: q<=8'h02;
	15'h17eb: q<=8'hc9;
	15'h17ec: q<=8'h10;
	15'h17ed: q<=8'hb0;
	15'h17ee: q<=8'h0c;
	15'h17ef: q<=8'hac;
	15'h17f0: q<=8'h15;
	15'h17f1: q<=8'h01;
	15'h17f2: q<=8'h10;
	15'h17f3: q<=8'h05;
	15'h17f4: q<=8'ha9;
	15'h17f5: q<=8'hf0;
	15'h17f6: q<=8'hb8;
	15'h17f7: q<=8'h50;
	15'h17f8: q<=8'h02;
	15'h17f9: q<=8'ha9;
	15'h17fa: q<=8'h00;
	15'h17fb: q<=8'hb8;
	15'h17fc: q<=8'h50;
	15'h17fd: q<=8'h20;
	15'h17fe: q<=8'hac;
	15'h17ff: q<=8'h15;
	15'h1800: q<=8'h01;
	15'h1801: q<=8'h10;
	15'h1802: q<=8'h1b;
	15'h1803: q<=8'h8a;
	15'h1804: q<=8'h18;
	15'h1805: q<=8'h69;
	15'h1806: q<=8'h01;
	15'h1807: q<=8'hc9;
	15'h1808: q<=8'h08;
	15'h1809: q<=8'h90;
	15'h180a: q<=8'h02;
	15'h180b: q<=8'ha9;
	15'h180c: q<=8'h00;
	15'h180d: q<=8'ha8;
	15'h180e: q<=8'hb9;
	15'h180f: q<=8'hfe;
	15'h1810: q<=8'h03;
	15'h1811: q<=8'hf0;
	15'h1812: q<=8'h0b;
	15'h1813: q<=8'hc9;
	15'h1814: q<=8'hd5;
	15'h1815: q<=8'hb0;
	15'h1816: q<=8'h05;
	15'h1817: q<=8'ha9;
	15'h1818: q<=8'hf0;
	15'h1819: q<=8'hb8;
	15'h181a: q<=8'h50;
	15'h181b: q<=8'h02;
	15'h181c: q<=8'ha9;
	15'h181d: q<=8'h00;
	15'h181e: q<=8'h9d;
	15'h181f: q<=8'hfe;
	15'h1820: q<=8'h03;
	15'h1821: q<=8'h05;
	15'h1822: q<=8'h29;
	15'h1823: q<=8'h85;
	15'h1824: q<=8'h29;
	15'h1825: q<=8'hc6;
	15'h1826: q<=8'h37;
	15'h1827: q<=8'h10;
	15'h1828: q<=8'hb6;
	15'h1829: q<=8'ha5;
	15'h182a: q<=8'h29;
	15'h182b: q<=8'hd0;
	15'h182c: q<=8'h03;
	15'h182d: q<=8'h8d;
	15'h182e: q<=8'h15;
	15'h182f: q<=8'h01;
	15'h1830: q<=8'h60;
	15'h1831: q<=8'ha9;
	15'h1832: q<=8'h00;
	15'h1833: q<=8'h8d;
	15'h1834: q<=8'haa;
	15'h1835: q<=8'h03;
	15'h1836: q<=8'h8d;
	15'h1837: q<=8'h25;
	15'h1838: q<=8'h01;
	15'h1839: q<=8'h60;
	15'h183a: q<=8'ha5;
	15'h183b: q<=8'h05;
	15'h183c: q<=8'h10;
	15'h183d: q<=8'h3e;
	15'h183e: q<=8'had;
	15'h183f: q<=8'h25;
	15'h1840: q<=8'h01;
	15'h1841: q<=8'hd0;
	15'h1842: q<=8'h23;
	15'h1843: q<=8'had;
	15'h1844: q<=8'h01;
	15'h1845: q<=8'h02;
	15'h1846: q<=8'h30;
	15'h1847: q<=8'h1b;
	15'h1848: q<=8'ha5;
	15'h1849: q<=8'h4e;
	15'h184a: q<=8'h29;
	15'h184b: q<=8'h08;
	15'h184c: q<=8'hf0;
	15'h184d: q<=8'h15;
	15'h184e: q<=8'had;
	15'h184f: q<=8'haa;
	15'h1850: q<=8'h03;
	15'h1851: q<=8'hc9;
	15'h1852: q<=8'h02;
	15'h1853: q<=8'hb0;
	15'h1854: q<=8'h08;
	15'h1855: q<=8'hee;
	15'h1856: q<=8'haa;
	15'h1857: q<=8'h03;
	15'h1858: q<=8'ha9;
	15'h1859: q<=8'h01;
	15'h185a: q<=8'h8d;
	15'h185b: q<=8'h25;
	15'h185c: q<=8'h01;
	15'h185d: q<=8'ha5;
	15'h185e: q<=8'h4e;
	15'h185f: q<=8'h29;
	15'h1860: q<=8'h77;
	15'h1861: q<=8'h85;
	15'h1862: q<=8'h4e;
	15'h1863: q<=8'hb8;
	15'h1864: q<=8'h50;
	15'h1865: q<=8'h16;
	15'h1866: q<=8'hee;
	15'h1867: q<=8'h25;
	15'h1868: q<=8'h01;
	15'h1869: q<=8'hae;
	15'h186a: q<=8'haa;
	15'h186b: q<=8'h03;
	15'h186c: q<=8'had;
	15'h186d: q<=8'h25;
	15'h186e: q<=8'h01;
	15'h186f: q<=8'hdd;
	15'h1870: q<=8'h83;
	15'h1871: q<=8'ha8;
	15'h1872: q<=8'h90;
	15'h1873: q<=8'h05;
	15'h1874: q<=8'ha9;
	15'h1875: q<=8'h00;
	15'h1876: q<=8'h8d;
	15'h1877: q<=8'h25;
	15'h1878: q<=8'h01;
	15'h1879: q<=8'h20;
	15'h187a: q<=8'h88;
	15'h187b: q<=8'ha8;
	15'h187c: q<=8'ha5;
	15'h187d: q<=8'h4e;
	15'h187e: q<=8'h29;
	15'h187f: q<=8'h7f;
	15'h1880: q<=8'h85;
	15'h1881: q<=8'h4e;
	15'h1882: q<=8'h60;
	15'h1883: q<=8'h00;
	15'h1884: q<=8'h13;
	15'h1885: q<=8'h05;
	15'h1886: q<=8'h00;
	15'h1887: q<=8'h00;
	15'h1888: q<=8'had;
	15'h1889: q<=8'h25;
	15'h188a: q<=8'h01;
	15'h188b: q<=8'hc9;
	15'h188c: q<=8'h03;
	15'h188d: q<=8'h90;
	15'h188e: q<=8'h14;
	15'h188f: q<=8'h29;
	15'h1890: q<=8'h01;
	15'h1891: q<=8'hd0;
	15'h1892: q<=8'h10;
	15'h1893: q<=8'hac;
	15'h1894: q<=8'h1c;
	15'h1895: q<=8'h01;
	15'h1896: q<=8'hb9;
	15'h1897: q<=8'hdf;
	15'h1898: q<=8'h02;
	15'h1899: q<=8'hd0;
	15'h189a: q<=8'h09;
	15'h189b: q<=8'h88;
	15'h189c: q<=8'h10;
	15'h189d: q<=8'hf8;
	15'h189e: q<=8'ha9;
	15'h189f: q<=8'h00;
	15'h18a0: q<=8'h8d;
	15'h18a1: q<=8'h25;
	15'h18a2: q<=8'h01;
	15'h18a3: q<=8'h60;
	15'h18a4: q<=8'hb9;
	15'h18a5: q<=8'h8a;
	15'h18a6: q<=8'h02;
	15'h18a7: q<=8'h29;
	15'h18a8: q<=8'hfc;
	15'h18a9: q<=8'h99;
	15'h18aa: q<=8'h8a;
	15'h18ab: q<=8'h02;
	15'h18ac: q<=8'h4c;
	15'h18ad: q<=8'h98;
	15'h18ae: q<=8'ha3;
	15'h18af: q<=8'he1;
	15'h18b0: q<=8'h24;
	15'h18b1: q<=8'h26;
	15'h18b2: q<=8'h28;
	15'h18b3: q<=8'h2a;
	15'h18b4: q<=8'ha9;
	15'h18b5: q<=8'h01;
	15'h18b6: q<=8'h85;
	15'h18b7: q<=8'h72;
	15'h18b8: q<=8'h20;
	15'h18b9: q<=8'h6a;
	15'h18ba: q<=8'hdf;
	15'h18bb: q<=8'ha0;
	15'h18bc: q<=8'h05;
	15'h18bd: q<=8'h20;
	15'h18be: q<=8'hd1;
	15'h18bf: q<=8'hb0;
	15'h18c0: q<=8'ha5;
	15'h18c1: q<=8'h05;
	15'h18c2: q<=8'h30;
	15'h18c3: q<=8'h26;
	15'h18c4: q<=8'ha2;
	15'h18c5: q<=8'h00;
	15'h18c6: q<=8'ha5;
	15'h18c7: q<=8'h03;
	15'h18c8: q<=8'h29;
	15'h18c9: q<=8'h20;
	15'h18ca: q<=8'hd0;
	15'h18cb: q<=8'h0c;
	15'h18cc: q<=8'ha2;
	15'h18cd: q<=8'h22;
	15'h18ce: q<=8'ha5;
	15'h18cf: q<=8'h06;
	15'h18d0: q<=8'hf0;
	15'h18d1: q<=8'h06;
	15'h18d2: q<=8'h24;
	15'h18d3: q<=8'ha2;
	15'h18d4: q<=8'h30;
	15'h18d5: q<=8'h02;
	15'h18d6: q<=8'ha2;
	15'h18d7: q<=8'h06;
	15'h18d8: q<=8'h20;
	15'h18d9: q<=8'h14;
	15'h18da: q<=8'hab;
	15'h18db: q<=8'h20;
	15'h18dc: q<=8'h0d;
	15'h18dd: q<=8'hab;
	15'h18de: q<=8'had;
	15'h18df: q<=8'he4;
	15'h18e0: q<=8'h31;
	15'h18e1: q<=8'h8d;
	15'h18e2: q<=8'ha6;
	15'h18e3: q<=8'h2f;
	15'h18e4: q<=8'h8d;
	15'h18e5: q<=8'ha8;
	15'h18e6: q<=8'h2f;
	15'h18e7: q<=8'h20;
	15'h18e8: q<=8'ha8;
	15'h18e9: q<=8'haa;
	15'h18ea: q<=8'ha9;
	15'h18eb: q<=8'h01;
	15'h18ec: q<=8'ha0;
	15'h18ed: q<=8'h00;
	15'h18ee: q<=8'h20;
	15'h18ef: q<=8'h7f;
	15'h18f0: q<=8'ha9;
	15'h18f1: q<=8'h24;
	15'h18f2: q<=8'h05;
	15'h18f3: q<=8'h30;
	15'h18f4: q<=8'h09;
	15'h18f5: q<=8'ha5;
	15'h18f6: q<=8'h43;
	15'h18f7: q<=8'h05;
	15'h18f8: q<=8'h44;
	15'h18f9: q<=8'h05;
	15'h18fa: q<=8'h45;
	15'h18fb: q<=8'hb8;
	15'h18fc: q<=8'h50;
	15'h18fd: q<=8'h02;
	15'h18fe: q<=8'ha5;
	15'h18ff: q<=8'h3e;
	15'h1900: q<=8'hf0;
	15'h1901: q<=8'h06;
	15'h1902: q<=8'ha9;
	15'h1903: q<=8'h01;
	15'h1904: q<=8'ha8;
	15'h1905: q<=8'h20;
	15'h1906: q<=8'h7f;
	15'h1907: q<=8'ha9;
	15'h1908: q<=8'ha5;
	15'h1909: q<=8'h00;
	15'h190a: q<=8'hc9;
	15'h190b: q<=8'h04;
	15'h190c: q<=8'hf0;
	15'h190d: q<=8'h35;
	15'h190e: q<=8'ha9;
	15'h190f: q<=8'h1d;
	15'h1910: q<=8'h85;
	15'h1911: q<=8'h3b;
	15'h1912: q<=8'ha9;
	15'h1913: q<=8'h07;
	15'h1914: q<=8'h85;
	15'h1915: q<=8'h3c;
	15'h1916: q<=8'hae;
	15'h1917: q<=8'he4;
	15'h1918: q<=8'hcd;
	15'h1919: q<=8'h20;
	15'h191a: q<=8'hd7;
	15'h191b: q<=8'ha9;
	15'h191c: q<=8'ha0;
	15'h191d: q<=8'h0a;
	15'h191e: q<=8'ha9;
	15'h191f: q<=8'ha7;
	15'h1920: q<=8'h59;
	15'h1921: q<=8'hce;
	15'h1922: q<=8'haa;
	15'h1923: q<=8'h88;
	15'h1924: q<=8'h10;
	15'h1925: q<=8'hfa;
	15'h1926: q<=8'h8d;
	15'h1927: q<=8'h6c;
	15'h1928: q<=8'h01;
	15'h1929: q<=8'hae;
	15'h192a: q<=8'he5;
	15'h192b: q<=8'hcd;
	15'h192c: q<=8'ha9;
	15'h192d: q<=8'h02;
	15'h192e: q<=8'h85;
	15'h192f: q<=8'h38;
	15'h1930: q<=8'ha4;
	15'h1931: q<=8'h38;
	15'h1932: q<=8'hb9;
	15'h1933: q<=8'h1b;
	15'h1934: q<=8'h06;
	15'h1935: q<=8'h0a;
	15'h1936: q<=8'ha8;
	15'h1937: q<=8'hb9;
	15'h1938: q<=8'hfa;
	15'h1939: q<=8'h31;
	15'h193a: q<=8'h9d;
	15'h193b: q<=8'h60;
	15'h193c: q<=8'h2f;
	15'h193d: q<=8'he8;
	15'h193e: q<=8'he8;
	15'h193f: q<=8'hc6;
	15'h1940: q<=8'h38;
	15'h1941: q<=8'h10;
	15'h1942: q<=8'hed;
	15'h1943: q<=8'ha9;
	15'h1944: q<=8'h2f;
	15'h1945: q<=8'ha2;
	15'h1946: q<=8'h60;
	15'h1947: q<=8'h20;
	15'h1948: q<=8'h39;
	15'h1949: q<=8'hdf;
	15'h194a: q<=8'had;
	15'h194b: q<=8'h23;
	15'h194c: q<=8'h01;
	15'h194d: q<=8'h10;
	15'h194e: q<=8'h05;
	15'h194f: q<=8'ha2;
	15'h1950: q<=8'h36;
	15'h1951: q<=8'h20;
	15'h1952: q<=8'h14;
	15'h1953: q<=8'hab;
	15'h1954: q<=8'ha5;
	15'h1955: q<=8'h00;
	15'h1956: q<=8'hc9;
	15'h1957: q<=8'h18;
	15'h1958: q<=8'hd0;
	15'h1959: q<=8'h22;
	15'h195a: q<=8'ha5;
	15'h195b: q<=8'h05;
	15'h195c: q<=8'h10;
	15'h195d: q<=8'h1e;
	15'h195e: q<=8'ha6;
	15'h195f: q<=8'h3d;
	15'h1960: q<=8'hbd;
	15'h1961: q<=8'h02;
	15'h1962: q<=8'h01;
	15'h1963: q<=8'hf0;
	15'h1964: q<=8'h0d;
	15'h1965: q<=8'ha2;
	15'h1966: q<=8'h30;
	15'h1967: q<=8'h20;
	15'h1968: q<=8'h14;
	15'h1969: q<=8'hab;
	15'h196a: q<=8'ha4;
	15'h196b: q<=8'h3d;
	15'h196c: q<=8'hbe;
	15'h196d: q<=8'h02;
	15'h196e: q<=8'h01;
	15'h196f: q<=8'h20;
	15'h1970: q<=8'hc6;
	15'h1971: q<=8'hb0;
	15'h1972: q<=8'ha2;
	15'h1973: q<=8'h3a;
	15'h1974: q<=8'h20;
	15'h1975: q<=8'h14;
	15'h1976: q<=8'hab;
	15'h1977: q<=8'ha2;
	15'h1978: q<=8'h38;
	15'h1979: q<=8'h20;
	15'h197a: q<=8'h14;
	15'h197b: q<=8'hab;
	15'h197c: q<=8'h60;
	15'h197d: q<=8'h42;
	15'h197e: q<=8'h45;
	15'h197f: q<=8'ha6;
	15'h1980: q<=8'h00;
	15'h1981: q<=8'he0;
	15'h1982: q<=8'h04;
	15'h1983: q<=8'h84;
	15'h1984: q<=8'h2b;
	15'h1985: q<=8'hc4;
	15'h1986: q<=8'h3d;
	15'h1987: q<=8'hd0;
	15'h1988: q<=8'h06;
	15'h1989: q<=8'h24;
	15'h198a: q<=8'h05;
	15'h198b: q<=8'h10;
	15'h198c: q<=8'h02;
	15'h198d: q<=8'ha9;
	15'h198e: q<=8'h00;
	15'h198f: q<=8'h09;
	15'h1990: q<=8'h70;
	15'h1991: q<=8'hbe;
	15'h1992: q<=8'hde;
	15'h1993: q<=8'hcd;
	15'h1994: q<=8'h9d;
	15'h1995: q<=8'h60;
	15'h1996: q<=8'h2f;
	15'h1997: q<=8'hbe;
	15'h1998: q<=8'he0;
	15'h1999: q<=8'hcd;
	15'h199a: q<=8'hb9;
	15'h199b: q<=8'h48;
	15'h199c: q<=8'h00;
	15'h199d: q<=8'h85;
	15'h199e: q<=8'h38;
	15'h199f: q<=8'hf0;
	15'h19a0: q<=8'h06;
	15'h19a1: q<=8'hc4;
	15'h19a2: q<=8'h3d;
	15'h19a3: q<=8'hd0;
	15'h19a4: q<=8'h02;
	15'h19a5: q<=8'hc6;
	15'h19a6: q<=8'h38;
	15'h19a7: q<=8'ha0;
	15'h19a8: q<=8'h01;
	15'h19a9: q<=8'had;
	15'h19aa: q<=8'h84;
	15'h19ab: q<=8'h32;
	15'h19ac: q<=8'hc4;
	15'h19ad: q<=8'h38;
	15'h19ae: q<=8'h90;
	15'h19af: q<=8'h05;
	15'h19b0: q<=8'hf0;
	15'h19b1: q<=8'h03;
	15'h19b2: q<=8'had;
	15'h19b3: q<=8'h86;
	15'h19b4: q<=8'h32;
	15'h19b5: q<=8'h9d;
	15'h19b6: q<=8'h60;
	15'h19b7: q<=8'h2f;
	15'h19b8: q<=8'he8;
	15'h19b9: q<=8'he8;
	15'h19ba: q<=8'hc8;
	15'h19bb: q<=8'hc0;
	15'h19bc: q<=8'h07;
	15'h19bd: q<=8'h90;
	15'h19be: q<=8'hea;
	15'h19bf: q<=8'ha4;
	15'h19c0: q<=8'h2b;
	15'h19c1: q<=8'ha5;
	15'h19c2: q<=8'h00;
	15'h19c3: q<=8'hc9;
	15'h19c4: q<=8'h04;
	15'h19c5: q<=8'hd0;
	15'h19c6: q<=8'h04;
	15'h19c7: q<=8'hc4;
	15'h19c8: q<=8'h3d;
	15'h19c9: q<=8'hd0;
	15'h19ca: q<=8'h30;
	15'h19cb: q<=8'hbe;
	15'h19cc: q<=8'he2;
	15'h19cd: q<=8'hcd;
	15'h19ce: q<=8'hb9;
	15'h19cf: q<=8'h7d;
	15'h19d0: q<=8'ha9;
	15'h19d1: q<=8'h85;
	15'h19d2: q<=8'h3b;
	15'h19d3: q<=8'ha9;
	15'h19d4: q<=8'h00;
	15'h19d5: q<=8'h85;
	15'h19d6: q<=8'h3c;
	15'h19d7: q<=8'ha0;
	15'h19d8: q<=8'h02;
	15'h19d9: q<=8'h84;
	15'h19da: q<=8'h2a;
	15'h19db: q<=8'h38;
	15'h19dc: q<=8'h08;
	15'h19dd: q<=8'ha0;
	15'h19de: q<=8'h00;
	15'h19df: q<=8'hb1;
	15'h19e0: q<=8'h3b;
	15'h19e1: q<=8'h4a;
	15'h19e2: q<=8'h4a;
	15'h19e3: q<=8'h4a;
	15'h19e4: q<=8'h4a;
	15'h19e5: q<=8'h28;
	15'h19e6: q<=8'h20;
	15'h19e7: q<=8'hfc;
	15'h19e8: q<=8'ha9;
	15'h19e9: q<=8'ha5;
	15'h19ea: q<=8'h2a;
	15'h19eb: q<=8'hd0;
	15'h19ec: q<=8'h01;
	15'h19ed: q<=8'h18;
	15'h19ee: q<=8'ha0;
	15'h19ef: q<=8'h00;
	15'h19f0: q<=8'hb1;
	15'h19f1: q<=8'h3b;
	15'h19f2: q<=8'h20;
	15'h19f3: q<=8'hfc;
	15'h19f4: q<=8'ha9;
	15'h19f5: q<=8'hc6;
	15'h19f6: q<=8'h3b;
	15'h19f7: q<=8'hc6;
	15'h19f8: q<=8'h2a;
	15'h19f9: q<=8'h10;
	15'h19fa: q<=8'he1;
	15'h19fb: q<=8'h60;
	15'h19fc: q<=8'h29;
	15'h19fd: q<=8'h0f;
	15'h19fe: q<=8'ha8;
	15'h19ff: q<=8'hf0;
	15'h1a00: q<=8'h01;
	15'h1a01: q<=8'h18;
	15'h1a02: q<=8'hb0;
	15'h1a03: q<=8'h01;
	15'h1a04: q<=8'hc8;
	15'h1a05: q<=8'h08;
	15'h1a06: q<=8'h98;
	15'h1a07: q<=8'h0a;
	15'h1a08: q<=8'ha8;
	15'h1a09: q<=8'hb9;
	15'h1a0a: q<=8'he4;
	15'h1a0b: q<=8'h31;
	15'h1a0c: q<=8'h9d;
	15'h1a0d: q<=8'h60;
	15'h1a0e: q<=8'h2f;
	15'h1a0f: q<=8'he8;
	15'h1a10: q<=8'he8;
	15'h1a11: q<=8'h28;
	15'h1a12: q<=8'h60;
	15'h1a13: q<=8'ha6;
	15'h1a14: q<=8'h3e;
	15'h1a15: q<=8'h24;
	15'h1a16: q<=8'h05;
	15'h1a17: q<=8'h30;
	15'h1a18: q<=8'h0a;
	15'h1a19: q<=8'ha5;
	15'h1a1a: q<=8'h43;
	15'h1a1b: q<=8'h05;
	15'h1a1c: q<=8'h44;
	15'h1a1d: q<=8'h05;
	15'h1a1e: q<=8'h45;
	15'h1a1f: q<=8'hf0;
	15'h1a20: q<=8'h02;
	15'h1a21: q<=8'ha2;
	15'h1a22: q<=8'h01;
	15'h1a23: q<=8'ha9;
	15'h1a24: q<=8'h60;
	15'h1a25: q<=8'h85;
	15'h1a26: q<=8'h74;
	15'h1a27: q<=8'ha9;
	15'h1a28: q<=8'h2f;
	15'h1a29: q<=8'h85;
	15'h1a2a: q<=8'h75;
	15'h1a2b: q<=8'hbd;
	15'h1a2c: q<=8'h66;
	15'h1a2d: q<=8'hce;
	15'h1a2e: q<=8'ha8;
	15'h1a2f: q<=8'h38;
	15'h1a30: q<=8'h65;
	15'h1a31: q<=8'h74;
	15'h1a32: q<=8'h48;
	15'h1a33: q<=8'hb9;
	15'h1a34: q<=8'he6;
	15'h1a35: q<=8'hcd;
	15'h1a36: q<=8'h91;
	15'h1a37: q<=8'h74;
	15'h1a38: q<=8'h88;
	15'h1a39: q<=8'hd0;
	15'h1a3a: q<=8'hf8;
	15'h1a3b: q<=8'hb9;
	15'h1a3c: q<=8'he6;
	15'h1a3d: q<=8'hcd;
	15'h1a3e: q<=8'h91;
	15'h1a3f: q<=8'h74;
	15'h1a40: q<=8'ha5;
	15'h1a41: q<=8'h05;
	15'h1a42: q<=8'h10;
	15'h1a43: q<=8'h10;
	15'h1a44: q<=8'ha9;
	15'h1a45: q<=8'h2f;
	15'h1a46: q<=8'h85;
	15'h1a47: q<=8'h75;
	15'h1a48: q<=8'ha9;
	15'h1a49: q<=8'ha6;
	15'h1a4a: q<=8'h85;
	15'h1a4b: q<=8'h74;
	15'h1a4c: q<=8'ha5;
	15'h1a4d: q<=8'h9f;
	15'h1a4e: q<=8'h18;
	15'h1a4f: q<=8'h69;
	15'h1a50: q<=8'h01;
	15'h1a51: q<=8'h20;
	15'h1a52: q<=8'h77;
	15'h1a53: q<=8'haf;
	15'h1a54: q<=8'h68;
	15'h1a55: q<=8'h85;
	15'h1a56: q<=8'h74;
	15'h1a57: q<=8'h4c;
	15'h1a58: q<=8'h09;
	15'h1a59: q<=8'hdf;
	15'h1a5a: q<=8'ha2;
	15'h1a5b: q<=8'h08;
	15'h1a5c: q<=8'h20;
	15'h1a5d: q<=8'h14;
	15'h1a5e: q<=8'hab;
	15'h1a5f: q<=8'h4c;
	15'h1a60: q<=8'h69;
	15'h1a61: q<=8'haa;
	15'h1a62: q<=8'ha9;
	15'h1a63: q<=8'h30;
	15'h1a64: q<=8'ha2;
	15'h1a65: q<=8'h00;
	15'h1a66: q<=8'h20;
	15'h1a67: q<=8'h17;
	15'h1a68: q<=8'hab;
	15'h1a69: q<=8'h20;
	15'h1a6a: q<=8'h92;
	15'h1a6b: q<=8'haa;
	15'h1a6c: q<=8'h4c;
	15'h1a6d: q<=8'he7;
	15'h1a6e: q<=8'ha8;
	15'h1a6f: q<=8'h20;
	15'h1a70: q<=8'hb4;
	15'h1a71: q<=8'ha8;
	15'h1a72: q<=8'ha9;
	15'h1a73: q<=8'h00;
	15'h1a74: q<=8'ha2;
	15'h1a75: q<=8'h06;
	15'h1a76: q<=8'h4c;
	15'h1a77: q<=8'h17;
	15'h1a78: q<=8'hab;
	15'h1a79: q<=8'ha9;
	15'h1a7a: q<=8'h00;
	15'h1a7b: q<=8'ha2;
	15'h1a7c: q<=8'h32;
	15'h1a7d: q<=8'h20;
	15'h1a7e: q<=8'h17;
	15'h1a7f: q<=8'hab;
	15'h1a80: q<=8'ha5;
	15'h1a81: q<=8'h03;
	15'h1a82: q<=8'h29;
	15'h1a83: q<=8'h1f;
	15'h1a84: q<=8'hc9;
	15'h1a85: q<=8'h10;
	15'h1a86: q<=8'hb0;
	15'h1a87: q<=8'h07;
	15'h1a88: q<=8'ha9;
	15'h1a89: q<=8'he0;
	15'h1a8a: q<=8'ha2;
	15'h1a8b: q<=8'h22;
	15'h1a8c: q<=8'h20;
	15'h1a8d: q<=8'h17;
	15'h1a8e: q<=8'hab;
	15'h1a8f: q<=8'h4c;
	15'h1a90: q<=8'hb4;
	15'h1a91: q<=8'ha8;
	15'h1a92: q<=8'ha2;
	15'h1a93: q<=8'h02;
	15'h1a94: q<=8'h20;
	15'h1a95: q<=8'h14;
	15'h1a96: q<=8'hab;
	15'h1a97: q<=8'ha9;
	15'h1a98: q<=8'h00;
	15'h1a99: q<=8'h20;
	15'h1a9a: q<=8'hdd;
	15'h1a9b: q<=8'hb0;
	15'h1a9c: q<=8'ha6;
	15'h1a9d: q<=8'h3d;
	15'h1a9e: q<=8'he8;
	15'h1a9f: q<=8'h86;
	15'h1aa0: q<=8'h61;
	15'h1aa1: q<=8'ha9;
	15'h1aa2: q<=8'h61;
	15'h1aa3: q<=8'ha0;
	15'h1aa4: q<=8'h01;
	15'h1aa5: q<=8'h4c;
	15'h1aa6: q<=8'hb1;
	15'h1aa7: q<=8'hdf;
	15'h1aa8: q<=8'ha5;
	15'h1aa9: q<=8'h09;
	15'h1aaa: q<=8'h29;
	15'h1aab: q<=8'h03;
	15'h1aac: q<=8'haa;
	15'h1aad: q<=8'hbd;
	15'h1aae: q<=8'hb0;
	15'h1aaf: q<=8'ha8;
	15'h1ab0: q<=8'haa;
	15'h1ab1: q<=8'h20;
	15'h1ab2: q<=8'h14;
	15'h1ab3: q<=8'hab;
	15'h1ab4: q<=8'hce;
	15'h1ab5: q<=8'h6e;
	15'h1ab6: q<=8'h01;
	15'h1ab7: q<=8'ha5;
	15'h1ab8: q<=8'h0a;
	15'h1ab9: q<=8'h29;
	15'h1aba: q<=8'h01;
	15'h1abb: q<=8'hf0;
	15'h1abc: q<=8'h0e;
	15'h1abd: q<=8'ha5;
	15'h1abe: q<=8'h03;
	15'h1abf: q<=8'h29;
	15'h1ac0: q<=8'h20;
	15'h1ac1: q<=8'hd0;
	15'h1ac2: q<=8'h08;
	15'h1ac3: q<=8'ha2;
	15'h1ac4: q<=8'h32;
	15'h1ac5: q<=8'h20;
	15'h1ac6: q<=8'h14;
	15'h1ac7: q<=8'hab;
	15'h1ac8: q<=8'hb8;
	15'h1ac9: q<=8'h50;
	15'h1aca: q<=8'h03;
	15'h1acb: q<=8'h20;
	15'h1acc: q<=8'hca;
	15'h1acd: q<=8'hae;
	15'h1ace: q<=8'ha2;
	15'h1acf: q<=8'h2c;
	15'h1ad0: q<=8'h20;
	15'h1ad1: q<=8'h14;
	15'h1ad2: q<=8'hab;
	15'h1ad3: q<=8'ha2;
	15'h1ad4: q<=8'h2e;
	15'h1ad5: q<=8'h20;
	15'h1ad6: q<=8'h14;
	15'h1ad7: q<=8'hab;
	15'h1ad8: q<=8'ha5;
	15'h1ad9: q<=8'h06;
	15'h1ada: q<=8'hc9;
	15'h1adb: q<=8'h28;
	15'h1adc: q<=8'h90;
	15'h1add: q<=8'h04;
	15'h1ade: q<=8'ha9;
	15'h1adf: q<=8'h28;
	15'h1ae0: q<=8'h85;
	15'h1ae1: q<=8'h06;
	15'h1ae2: q<=8'h20;
	15'h1ae3: q<=8'h77;
	15'h1ae4: q<=8'haf;
	15'h1ae5: q<=8'ha5;
	15'h1ae6: q<=8'h17;
	15'h1ae7: q<=8'hf0;
	15'h1ae8: q<=8'h09;
	15'h1ae9: q<=8'had;
	15'h1aea: q<=8'hf4;
	15'h1aeb: q<=8'haa;
	15'h1aec: q<=8'hae;
	15'h1aed: q<=8'hf3;
	15'h1aee: q<=8'haa;
	15'h1aef: q<=8'h20;
	15'h1af0: q<=8'h39;
	15'h1af1: q<=8'hdf;
	15'h1af2: q<=8'h60;
	15'h1af3: q<=8'h5c;
	15'h1af4: q<=8'h32;
	15'h1af5: q<=8'hf8;
	15'h1af6: q<=8'h85;
	15'h1af7: q<=8'h29;
	15'h1af8: q<=8'ha9;
	15'h1af9: q<=8'h00;
	15'h1afa: q<=8'h85;
	15'h1afb: q<=8'h2c;
	15'h1afc: q<=8'ha0;
	15'h1afd: q<=8'h07;
	15'h1afe: q<=8'h06;
	15'h1aff: q<=8'h29;
	15'h1b00: q<=8'ha5;
	15'h1b01: q<=8'h2c;
	15'h1b02: q<=8'h65;
	15'h1b03: q<=8'h2c;
	15'h1b04: q<=8'h85;
	15'h1b05: q<=8'h2c;
	15'h1b06: q<=8'h88;
	15'h1b07: q<=8'h10;
	15'h1b08: q<=8'hf5;
	15'h1b09: q<=8'hd8;
	15'h1b0a: q<=8'h85;
	15'h1b0b: q<=8'h29;
	15'h1b0c: q<=8'h60;
	15'h1b0d: q<=8'ha9;
	15'h1b0e: q<=8'h20;
	15'h1b0f: q<=8'ha2;
	15'h1b10: q<=8'h80;
	15'h1b11: q<=8'h4c;
	15'h1b12: q<=8'h57;
	15'h1b13: q<=8'hdf;
	15'h1b14: q<=8'hbd;
	15'h1b15: q<=8'h22;
	15'h1b16: q<=8'hd1;
	15'h1b17: q<=8'h86;
	15'h1b18: q<=8'h35;
	15'h1b19: q<=8'h85;
	15'h1b1a: q<=8'h2b;
	15'h1b1b: q<=8'ha4;
	15'h1b1c: q<=8'h35;
	15'h1b1d: q<=8'hb1;
	15'h1b1e: q<=8'hac;
	15'h1b1f: q<=8'h85;
	15'h1b20: q<=8'h3b;
	15'h1b21: q<=8'hc8;
	15'h1b22: q<=8'hb1;
	15'h1b23: q<=8'hac;
	15'h1b24: q<=8'h85;
	15'h1b25: q<=8'h3c;
	15'h1b26: q<=8'he0;
	15'h1b27: q<=8'h2c;
	15'h1b28: q<=8'hd0;
	15'h1b29: q<=8'h08;
	15'h1b2a: q<=8'ha5;
	15'h1b2b: q<=8'h74;
	15'h1b2c: q<=8'h85;
	15'h1b2d: q<=8'hb6;
	15'h1b2e: q<=8'ha5;
	15'h1b2f: q<=8'h75;
	15'h1b30: q<=8'h85;
	15'h1b31: q<=8'hb7;
	15'h1b32: q<=8'ha0;
	15'h1b33: q<=8'h00;
	15'h1b34: q<=8'hb1;
	15'h1b35: q<=8'h3b;
	15'h1b36: q<=8'h85;
	15'h1b37: q<=8'h2a;
	15'h1b38: q<=8'h20;
	15'h1b39: q<=8'h0d;
	15'h1b3a: q<=8'hab;
	15'h1b3b: q<=8'ha9;
	15'h1b3c: q<=8'h00;
	15'h1b3d: q<=8'h85;
	15'h1b3e: q<=8'h73;
	15'h1b3f: q<=8'ha9;
	15'h1b40: q<=8'h01;
	15'h1b41: q<=8'h85;
	15'h1b42: q<=8'h72;
	15'h1b43: q<=8'h20;
	15'h1b44: q<=8'h6a;
	15'h1b45: q<=8'hdf;
	15'h1b46: q<=8'ha5;
	15'h1b47: q<=8'h2a;
	15'h1b48: q<=8'ha6;
	15'h1b49: q<=8'h2b;
	15'h1b4a: q<=8'h20;
	15'h1b4b: q<=8'h75;
	15'h1b4c: q<=8'hdf;
	15'h1b4d: q<=8'ha4;
	15'h1b4e: q<=8'h35;
	15'h1b4f: q<=8'hb1;
	15'h1b50: q<=8'hac;
	15'h1b51: q<=8'h85;
	15'h1b52: q<=8'h3b;
	15'h1b53: q<=8'hc8;
	15'h1b54: q<=8'hb1;
	15'h1b55: q<=8'hac;
	15'h1b56: q<=8'h85;
	15'h1b57: q<=8'h3c;
	15'h1b58: q<=8'ha6;
	15'h1b59: q<=8'h35;
	15'h1b5a: q<=8'hbd;
	15'h1b5b: q<=8'h21;
	15'h1b5c: q<=8'hd1;
	15'h1b5d: q<=8'h48;
	15'h1b5e: q<=8'h4a;
	15'h1b5f: q<=8'h4a;
	15'h1b60: q<=8'h4a;
	15'h1b61: q<=8'h4a;
	15'h1b62: q<=8'ha8;
	15'h1b63: q<=8'h20;
	15'h1b64: q<=8'hd1;
	15'h1b65: q<=8'hb0;
	15'h1b66: q<=8'h68;
	15'h1b67: q<=8'h29;
	15'h1b68: q<=8'h0f;
	15'h1b69: q<=8'h20;
	15'h1b6a: q<=8'hdd;
	15'h1b6b: q<=8'hb0;
	15'h1b6c: q<=8'ha0;
	15'h1b6d: q<=8'h01;
	15'h1b6e: q<=8'ha9;
	15'h1b6f: q<=8'h00;
	15'h1b70: q<=8'h85;
	15'h1b71: q<=8'h2a;
	15'h1b72: q<=8'hb1;
	15'h1b73: q<=8'h3b;
	15'h1b74: q<=8'h85;
	15'h1b75: q<=8'h2b;
	15'h1b76: q<=8'h29;
	15'h1b77: q<=8'h7f;
	15'h1b78: q<=8'hc8;
	15'h1b79: q<=8'h84;
	15'h1b7a: q<=8'h2c;
	15'h1b7b: q<=8'haa;
	15'h1b7c: q<=8'hbd;
	15'h1b7d: q<=8'he4;
	15'h1b7e: q<=8'h31;
	15'h1b7f: q<=8'ha4;
	15'h1b80: q<=8'h2a;
	15'h1b81: q<=8'h91;
	15'h1b82: q<=8'h74;
	15'h1b83: q<=8'hc8;
	15'h1b84: q<=8'hbd;
	15'h1b85: q<=8'he5;
	15'h1b86: q<=8'h31;
	15'h1b87: q<=8'h91;
	15'h1b88: q<=8'h74;
	15'h1b89: q<=8'hc8;
	15'h1b8a: q<=8'h84;
	15'h1b8b: q<=8'h2a;
	15'h1b8c: q<=8'ha4;
	15'h1b8d: q<=8'h2c;
	15'h1b8e: q<=8'h24;
	15'h1b8f: q<=8'h2b;
	15'h1b90: q<=8'h10;
	15'h1b91: q<=8'he0;
	15'h1b92: q<=8'ha4;
	15'h1b93: q<=8'h2a;
	15'h1b94: q<=8'h88;
	15'h1b95: q<=8'h4c;
	15'h1b96: q<=8'h5f;
	15'h1b97: q<=8'hdf;
	15'h1b98: q<=8'h86;
	15'h1b99: q<=8'h35;
	15'h1b9a: q<=8'h85;
	15'h1b9b: q<=8'h2a;
	15'h1b9c: q<=8'ha9;
	15'h1b9d: q<=8'h00;
	15'h1b9e: q<=8'h85;
	15'h1b9f: q<=8'h2b;
	15'h1ba0: q<=8'hf0;
	15'h1ba1: q<=8'h99;
	15'h1ba2: q<=8'h20;
	15'h1ba3: q<=8'h20;
	15'h1ba4: q<=8'hac;
	15'h1ba5: q<=8'had;
	15'h1ba6: q<=8'hc9;
	15'h1ba7: q<=8'h01;
	15'h1ba8: q<=8'h29;
	15'h1ba9: q<=8'h03;
	15'h1baa: q<=8'hf0;
	15'h1bab: q<=8'h5b;
	15'h1bac: q<=8'h20;
	15'h1bad: q<=8'h20;
	15'h1bae: q<=8'hac;
	15'h1baf: q<=8'ha9;
	15'h1bb0: q<=8'h08;
	15'h1bb1: q<=8'h8d;
	15'h1bb2: q<=8'h00;
	15'h1bb3: q<=8'h01;
	15'h1bb4: q<=8'had;
	15'h1bb5: q<=8'h1b;
	15'h1bb6: q<=8'h07;
	15'h1bb7: q<=8'h0d;
	15'h1bb8: q<=8'h1c;
	15'h1bb9: q<=8'h07;
	15'h1bba: q<=8'h0d;
	15'h1bbb: q<=8'h1d;
	15'h1bbc: q<=8'h07;
	15'h1bbd: q<=8'hd0;
	15'h1bbe: q<=8'h03;
	15'h1bbf: q<=8'h20;
	15'h1bc0: q<=8'h36;
	15'h1bc1: q<=8'hac;
	15'h1bc2: q<=8'ha2;
	15'h1bc3: q<=8'h17;
	15'h1bc4: q<=8'had;
	15'h1bc5: q<=8'hc9;
	15'h1bc6: q<=8'h01;
	15'h1bc7: q<=8'h29;
	15'h1bc8: q<=8'h01;
	15'h1bc9: q<=8'hd0;
	15'h1bca: q<=8'h02;
	15'h1bcb: q<=8'ha2;
	15'h1bcc: q<=8'h0e;
	15'h1bcd: q<=8'hbd;
	15'h1bce: q<=8'h08;
	15'h1bcf: q<=8'hac;
	15'h1bd0: q<=8'h9d;
	15'h1bd1: q<=8'h06;
	15'h1bd2: q<=8'h06;
	15'h1bd3: q<=8'hca;
	15'h1bd4: q<=8'h10;
	15'h1bd5: q<=8'hf7;
	15'h1bd6: q<=8'ha2;
	15'h1bd7: q<=8'h17;
	15'h1bd8: q<=8'had;
	15'h1bd9: q<=8'hc9;
	15'h1bda: q<=8'h01;
	15'h1bdb: q<=8'h29;
	15'h1bdc: q<=8'h02;
	15'h1bdd: q<=8'hd0;
	15'h1bde: q<=8'h02;
	15'h1bdf: q<=8'ha2;
	15'h1be0: q<=8'h0e;
	15'h1be1: q<=8'ha9;
	15'h1be2: q<=8'h01;
	15'h1be3: q<=8'h9d;
	15'h1be4: q<=8'h06;
	15'h1be5: q<=8'h07;
	15'h1be6: q<=8'hca;
	15'h1be7: q<=8'h10;
	15'h1be8: q<=8'hf8;
	15'h1be9: q<=8'had;
	15'h1bea: q<=8'hc9;
	15'h1beb: q<=8'h01;
	15'h1bec: q<=8'h29;
	15'h1bed: q<=8'h03;
	15'h1bee: q<=8'hf0;
	15'h1bef: q<=8'h0f;
	15'h1bf0: q<=8'ha5;
	15'h1bf1: q<=8'h0a;
	15'h1bf2: q<=8'h29;
	15'h1bf3: q<=8'hf8;
	15'h1bf4: q<=8'h8d;
	15'h1bf5: q<=8'h1e;
	15'h1bf6: q<=8'h07;
	15'h1bf7: q<=8'had;
	15'h1bf8: q<=8'h6a;
	15'h1bf9: q<=8'h01;
	15'h1bfa: q<=8'h29;
	15'h1bfb: q<=8'h03;
	15'h1bfc: q<=8'h8d;
	15'h1bfd: q<=8'h1f;
	15'h1bfe: q<=8'h07;
	15'h1bff: q<=8'had;
	15'h1c00: q<=8'hc9;
	15'h1c01: q<=8'h01;
	15'h1c02: q<=8'h29;
	15'h1c03: q<=8'hfc;
	15'h1c04: q<=8'h8d;
	15'h1c05: q<=8'hc9;
	15'h1c06: q<=8'h01;
	15'h1c07: q<=8'h60;
	15'h1c08: q<=8'h07;
	15'h1c09: q<=8'h04;
	15'h1c0a: q<=8'h01;
	15'h1c0b: q<=8'h0f;
	15'h1c0c: q<=8'h09;
	15'h1c0d: q<=8'h0c;
	15'h1c0e: q<=8'h0b;
	15'h1c0f: q<=8'h03;
	15'h1c10: q<=8'h12;
	15'h1c11: q<=8'h13;
	15'h1c12: q<=8'h05;
	15'h1c13: q<=8'h03;
	15'h1c14: q<=8'h07;
	15'h1c15: q<=8'h0f;
	15'h1c16: q<=8'h0c;
	15'h1c17: q<=8'h11;
	15'h1c18: q<=8'h11;
	15'h1c19: q<=8'h11;
	15'h1c1a: q<=8'h12;
	15'h1c1b: q<=8'h04;
	15'h1c1c: q<=8'h03;
	15'h1c1d: q<=8'h03;
	15'h1c1e: q<=8'h09;
	15'h1c1f: q<=8'h04;
	15'h1c20: q<=8'h20;
	15'h1c21: q<=8'hbb;
	15'h1c22: q<=8'hd6;
	15'h1c23: q<=8'ha5;
	15'h1c24: q<=8'h0a;
	15'h1c25: q<=8'h29;
	15'h1c26: q<=8'hf8;
	15'h1c27: q<=8'hcd;
	15'h1c28: q<=8'h1e;
	15'h1c29: q<=8'h07;
	15'h1c2a: q<=8'hd0;
	15'h1c2b: q<=8'h08;
	15'h1c2c: q<=8'had;
	15'h1c2d: q<=8'h6a;
	15'h1c2e: q<=8'h01;
	15'h1c2f: q<=8'h29;
	15'h1c30: q<=8'h03;
	15'h1c31: q<=8'hcd;
	15'h1c32: q<=8'h1f;
	15'h1c33: q<=8'h07;
	15'h1c34: q<=8'hf0;
	15'h1c35: q<=8'h08;
	15'h1c36: q<=8'had;
	15'h1c37: q<=8'hc9;
	15'h1c38: q<=8'h01;
	15'h1c39: q<=8'h09;
	15'h1c3a: q<=8'h03;
	15'h1c3b: q<=8'h8d;
	15'h1c3c: q<=8'hc9;
	15'h1c3d: q<=8'h01;
	15'h1c3e: q<=8'h60;
	15'h1c3f: q<=8'ha5;
	15'h1c40: q<=8'h05;
	15'h1c41: q<=8'h29;
	15'h1c42: q<=8'hbf;
	15'h1c43: q<=8'h85;
	15'h1c44: q<=8'h05;
	15'h1c45: q<=8'ha5;
	15'h1c46: q<=8'h09;
	15'h1c47: q<=8'h29;
	15'h1c48: q<=8'h43;
	15'h1c49: q<=8'hc9;
	15'h1c4a: q<=8'h40;
	15'h1c4b: q<=8'hd0;
	15'h1c4c: q<=8'h03;
	15'h1c4d: q<=8'h20;
	15'h1c4e: q<=8'h62;
	15'h1c4f: q<=8'hca;
	15'h1c50: q<=8'h20;
	15'h1c51: q<=8'hfb;
	15'h1c52: q<=8'hdd;
	15'h1c53: q<=8'ha9;
	15'h1c54: q<=8'h00;
	15'h1c55: q<=8'h8d;
	15'h1c56: q<=8'h01;
	15'h1c57: q<=8'h06;
	15'h1c58: q<=8'ha6;
	15'h1c59: q<=8'h3e;
	15'h1c5a: q<=8'hf0;
	15'h1c5b: q<=8'h02;
	15'h1c5c: q<=8'ha2;
	15'h1c5d: q<=8'h03;
	15'h1c5e: q<=8'hb5;
	15'h1c5f: q<=8'h42;
	15'h1c60: q<=8'h85;
	15'h1c61: q<=8'h2c;
	15'h1c62: q<=8'hb5;
	15'h1c63: q<=8'h41;
	15'h1c64: q<=8'h85;
	15'h1c65: q<=8'h2d;
	15'h1c66: q<=8'hb5;
	15'h1c67: q<=8'h40;
	15'h1c68: q<=8'h85;
	15'h1c69: q<=8'h2e;
	15'h1c6a: q<=8'h8a;
	15'h1c6b: q<=8'h29;
	15'h1c6c: q<=8'h01;
	15'h1c6d: q<=8'h85;
	15'h1c6e: q<=8'h36;
	15'h1c6f: q<=8'ha9;
	15'h1c70: q<=8'h00;
	15'h1c71: q<=8'h85;
	15'h1c72: q<=8'h2b;
	15'h1c73: q<=8'ha9;
	15'h1c74: q<=8'h1a;
	15'h1c75: q<=8'h85;
	15'h1c76: q<=8'h2a;
	15'h1c77: q<=8'h85;
	15'h1c78: q<=8'h29;
	15'h1c79: q<=8'ha9;
	15'h1c7a: q<=8'h00;
	15'h1c7b: q<=8'h8d;
	15'h1c7c: q<=8'h05;
	15'h1c7d: q<=8'h06;
	15'h1c7e: q<=8'ha0;
	15'h1c7f: q<=8'hfd;
	15'h1c80: q<=8'hb9;
	15'h1c81: q<=8'h20;
	15'h1c82: q<=8'h06;
	15'h1c83: q<=8'hc5;
	15'h1c84: q<=8'h2c;
	15'h1c85: q<=8'hd0;
	15'h1c86: q<=8'h14;
	15'h1c87: q<=8'hb9;
	15'h1c88: q<=8'h1f;
	15'h1c89: q<=8'h06;
	15'h1c8a: q<=8'hc5;
	15'h1c8b: q<=8'h2d;
	15'h1c8c: q<=8'hd0;
	15'h1c8d: q<=8'h0d;
	15'h1c8e: q<=8'hc0;
	15'h1c8f: q<=8'h52;
	15'h1c90: q<=8'h90;
	15'h1c91: q<=8'h08;
	15'h1c92: q<=8'hb9;
	15'h1c93: q<=8'h1e;
	15'h1c94: q<=8'h06;
	15'h1c95: q<=8'hc5;
	15'h1c96: q<=8'h2e;
	15'h1c97: q<=8'hb8;
	15'h1c98: q<=8'h50;
	15'h1c99: q<=8'h01;
	15'h1c9a: q<=8'h38;
	15'h1c9b: q<=8'hb0;
	15'h1c9c: q<=8'h4f;
	15'h1c9d: q<=8'hc0;
	15'h1c9e: q<=8'he8;
	15'h1c9f: q<=8'h90;
	15'h1ca0: q<=8'h1e;
	15'h1ca1: q<=8'ha5;
	15'h1ca2: q<=8'h29;
	15'h1ca3: q<=8'hbe;
	15'h1ca4: q<=8'h1e;
	15'h1ca5: q<=8'h05;
	15'h1ca6: q<=8'h99;
	15'h1ca7: q<=8'h1e;
	15'h1ca8: q<=8'h05;
	15'h1ca9: q<=8'h86;
	15'h1caa: q<=8'h29;
	15'h1cab: q<=8'ha5;
	15'h1cac: q<=8'h2a;
	15'h1cad: q<=8'hbe;
	15'h1cae: q<=8'h1f;
	15'h1caf: q<=8'h05;
	15'h1cb0: q<=8'h99;
	15'h1cb1: q<=8'h1f;
	15'h1cb2: q<=8'h05;
	15'h1cb3: q<=8'h86;
	15'h1cb4: q<=8'h2a;
	15'h1cb5: q<=8'ha5;
	15'h1cb6: q<=8'h2b;
	15'h1cb7: q<=8'hbe;
	15'h1cb8: q<=8'h20;
	15'h1cb9: q<=8'h05;
	15'h1cba: q<=8'h99;
	15'h1cbb: q<=8'h20;
	15'h1cbc: q<=8'h05;
	15'h1cbd: q<=8'h86;
	15'h1cbe: q<=8'h2b;
	15'h1cbf: q<=8'ha5;
	15'h1cc0: q<=8'h2d;
	15'h1cc1: q<=8'hbe;
	15'h1cc2: q<=8'h1f;
	15'h1cc3: q<=8'h06;
	15'h1cc4: q<=8'h99;
	15'h1cc5: q<=8'h1f;
	15'h1cc6: q<=8'h06;
	15'h1cc7: q<=8'h86;
	15'h1cc8: q<=8'h2d;
	15'h1cc9: q<=8'ha5;
	15'h1cca: q<=8'h2c;
	15'h1ccb: q<=8'hbe;
	15'h1ccc: q<=8'h20;
	15'h1ccd: q<=8'h06;
	15'h1cce: q<=8'h99;
	15'h1ccf: q<=8'h20;
	15'h1cd0: q<=8'h06;
	15'h1cd1: q<=8'h86;
	15'h1cd2: q<=8'h2c;
	15'h1cd3: q<=8'hc0;
	15'h1cd4: q<=8'h52;
	15'h1cd5: q<=8'h90;
	15'h1cd6: q<=8'h0a;
	15'h1cd7: q<=8'ha5;
	15'h1cd8: q<=8'h2e;
	15'h1cd9: q<=8'hbe;
	15'h1cda: q<=8'h1e;
	15'h1cdb: q<=8'h06;
	15'h1cdc: q<=8'h99;
	15'h1cdd: q<=8'h1e;
	15'h1cde: q<=8'h06;
	15'h1cdf: q<=8'h86;
	15'h1ce0: q<=8'h2e;
	15'h1ce1: q<=8'hc0;
	15'h1ce2: q<=8'h55;
	15'h1ce3: q<=8'h90;
	15'h1ce4: q<=8'h01;
	15'h1ce5: q<=8'h88;
	15'h1ce6: q<=8'h88;
	15'h1ce7: q<=8'h88;
	15'h1ce8: q<=8'hd0;
	15'h1ce9: q<=8'hb3;
	15'h1cea: q<=8'ha0;
	15'h1ceb: q<=8'h02;
	15'h1cec: q<=8'hee;
	15'h1ced: q<=8'h05;
	15'h1cee: q<=8'h06;
	15'h1cef: q<=8'hc0;
	15'h1cf0: q<=8'h55;
	15'h1cf1: q<=8'h90;
	15'h1cf2: q<=8'h01;
	15'h1cf3: q<=8'h88;
	15'h1cf4: q<=8'h88;
	15'h1cf5: q<=8'h88;
	15'h1cf6: q<=8'hd0;
	15'h1cf7: q<=8'h88;
	15'h1cf8: q<=8'ha6;
	15'h1cf9: q<=8'h36;
	15'h1cfa: q<=8'had;
	15'h1cfb: q<=8'h05;
	15'h1cfc: q<=8'h06;
	15'h1cfd: q<=8'h9d;
	15'h1cfe: q<=8'h00;
	15'h1cff: q<=8'h06;
	15'h1d00: q<=8'hca;
	15'h1d01: q<=8'h30;
	15'h1d02: q<=8'h03;
	15'h1d03: q<=8'h4c;
	15'h1d04: q<=8'h5e;
	15'h1d05: q<=8'hac;
	15'h1d06: q<=8'had;
	15'h1d07: q<=8'h01;
	15'h1d08: q<=8'h06;
	15'h1d09: q<=8'hcd;
	15'h1d0a: q<=8'h00;
	15'h1d0b: q<=8'h06;
	15'h1d0c: q<=8'h90;
	15'h1d0d: q<=8'h07;
	15'h1d0e: q<=8'hc9;
	15'h1d0f: q<=8'h63;
	15'h1d10: q<=8'hb0;
	15'h1d11: q<=8'h03;
	15'h1d12: q<=8'hee;
	15'h1d13: q<=8'h01;
	15'h1d14: q<=8'h06;
	15'h1d15: q<=8'ha5;
	15'h1d16: q<=8'h3d;
	15'h1d17: q<=8'h49;
	15'h1d18: q<=8'h01;
	15'h1d19: q<=8'h0a;
	15'h1d1a: q<=8'h0a;
	15'h1d1b: q<=8'h05;
	15'h1d1c: q<=8'h3d;
	15'h1d1d: q<=8'h69;
	15'h1d1e: q<=8'h05;
	15'h1d1f: q<=8'h8d;
	15'h1d20: q<=8'h03;
	15'h1d21: q<=8'h06;
	15'h1d22: q<=8'ha0;
	15'h1d23: q<=8'h14;
	15'h1d24: q<=8'had;
	15'h1d25: q<=8'h03;
	15'h1d26: q<=8'h06;
	15'h1d27: q<=8'hf0;
	15'h1d28: q<=8'h42;
	15'h1d29: q<=8'h29;
	15'h1d2a: q<=8'h03;
	15'h1d2b: q<=8'h85;
	15'h1d2c: q<=8'h3d;
	15'h1d2d: q<=8'hc6;
	15'h1d2e: q<=8'h3d;
	15'h1d2f: q<=8'h4e;
	15'h1d30: q<=8'h03;
	15'h1d31: q<=8'h06;
	15'h1d32: q<=8'h4e;
	15'h1d33: q<=8'h03;
	15'h1d34: q<=8'h06;
	15'h1d35: q<=8'ha6;
	15'h1d36: q<=8'h3d;
	15'h1d37: q<=8'hbd;
	15'h1d38: q<=8'h00;
	15'h1d39: q<=8'h06;
	15'h1d3a: q<=8'hf0;
	15'h1d3b: q<=8'h2c;
	15'h1d3c: q<=8'hc9;
	15'h1d3d: q<=8'h09;
	15'h1d3e: q<=8'hb0;
	15'h1d3f: q<=8'h28;
	15'h1d40: q<=8'h0a;
	15'h1d41: q<=8'h18;
	15'h1d42: q<=8'h7d;
	15'h1d43: q<=8'h00;
	15'h1d44: q<=8'h06;
	15'h1d45: q<=8'h49;
	15'h1d46: q<=8'hff;
	15'h1d47: q<=8'h38;
	15'h1d48: q<=8'he9;
	15'h1d49: q<=8'he5;
	15'h1d4a: q<=8'h8d;
	15'h1d4b: q<=8'h02;
	15'h1d4c: q<=8'h06;
	15'h1d4d: q<=8'h20;
	15'h1d4e: q<=8'h48;
	15'h1d4f: q<=8'hca;
	15'h1d50: q<=8'ha9;
	15'h1d51: q<=8'h60;
	15'h1d52: q<=8'h8d;
	15'h1d53: q<=8'h05;
	15'h1d54: q<=8'h06;
	15'h1d55: q<=8'ha9;
	15'h1d56: q<=8'h00;
	15'h1d57: q<=8'h85;
	15'h1d58: q<=8'h4e;
	15'h1d59: q<=8'h85;
	15'h1d5a: q<=8'h50;
	15'h1d5b: q<=8'ha9;
	15'h1d5c: q<=8'h02;
	15'h1d5d: q<=8'h8d;
	15'h1d5e: q<=8'h04;
	15'h1d5f: q<=8'h06;
	15'h1d60: q<=8'h20;
	15'h1d61: q<=8'h89;
	15'h1d62: q<=8'ha7;
	15'h1d63: q<=8'ha0;
	15'h1d64: q<=8'h24;
	15'h1d65: q<=8'h84;
	15'h1d66: q<=8'h00;
	15'h1d67: q<=8'h60;
	15'h1d68: q<=8'h4c;
	15'h1d69: q<=8'h22;
	15'h1d6a: q<=8'had;
	15'h1d6b: q<=8'h84;
	15'h1d6c: q<=8'h00;
	15'h1d6d: q<=8'h60;
	15'h1d6e: q<=8'ha9;
	15'h1d6f: q<=8'h06;
	15'h1d70: q<=8'h85;
	15'h1d71: q<=8'h01;
	15'h1d72: q<=8'ha5;
	15'h1d73: q<=8'h03;
	15'h1d74: q<=8'h29;
	15'h1d75: q<=8'h1f;
	15'h1d76: q<=8'hd0;
	15'h1d77: q<=8'h0a;
	15'h1d78: q<=8'hce;
	15'h1d79: q<=8'h05;
	15'h1d7a: q<=8'h06;
	15'h1d7b: q<=8'hd0;
	15'h1d7c: q<=8'h05;
	15'h1d7d: q<=8'ha0;
	15'h1d7e: q<=8'h14;
	15'h1d7f: q<=8'h84;
	15'h1d80: q<=8'h00;
	15'h1d81: q<=8'h60;
	15'h1d82: q<=8'hae;
	15'h1d83: q<=8'h02;
	15'h1d84: q<=8'h06;
	15'h1d85: q<=8'hbd;
	15'h1d86: q<=8'h06;
	15'h1d87: q<=8'h06;
	15'h1d88: q<=8'h20;
	15'h1d89: q<=8'hce;
	15'h1d8a: q<=8'had;
	15'h1d8b: q<=8'ha8;
	15'h1d8c: q<=8'h10;
	15'h1d8d: q<=8'h05;
	15'h1d8e: q<=8'ha9;
	15'h1d8f: q<=8'h1a;
	15'h1d90: q<=8'hb8;
	15'h1d91: q<=8'h50;
	15'h1d92: q<=8'h06;
	15'h1d93: q<=8'hc9;
	15'h1d94: q<=8'h1b;
	15'h1d95: q<=8'h90;
	15'h1d96: q<=8'h02;
	15'h1d97: q<=8'ha9;
	15'h1d98: q<=8'h00;
	15'h1d99: q<=8'hae;
	15'h1d9a: q<=8'h02;
	15'h1d9b: q<=8'h06;
	15'h1d9c: q<=8'h9d;
	15'h1d9d: q<=8'h06;
	15'h1d9e: q<=8'h06;
	15'h1d9f: q<=8'ha5;
	15'h1da0: q<=8'h4e;
	15'h1da1: q<=8'h29;
	15'h1da2: q<=8'h18;
	15'h1da3: q<=8'ha8;
	15'h1da4: q<=8'ha5;
	15'h1da5: q<=8'h4e;
	15'h1da6: q<=8'h29;
	15'h1da7: q<=8'h67;
	15'h1da8: q<=8'h85;
	15'h1da9: q<=8'h4e;
	15'h1daa: q<=8'h98;
	15'h1dab: q<=8'hf0;
	15'h1dac: q<=8'h20;
	15'h1dad: q<=8'hce;
	15'h1dae: q<=8'h02;
	15'h1daf: q<=8'h06;
	15'h1db0: q<=8'hce;
	15'h1db1: q<=8'h04;
	15'h1db2: q<=8'h06;
	15'h1db3: q<=8'h10;
	15'h1db4: q<=8'h12;
	15'h1db5: q<=8'ha6;
	15'h1db6: q<=8'h3d;
	15'h1db7: q<=8'hbd;
	15'h1db8: q<=8'h00;
	15'h1db9: q<=8'h06;
	15'h1dba: q<=8'hc9;
	15'h1dbb: q<=8'h04;
	15'h1dbc: q<=8'hb0;
	15'h1dbd: q<=8'h03;
	15'h1dbe: q<=8'h20;
	15'h1dbf: q<=8'hf7;
	15'h1dc0: q<=8'hdd;
	15'h1dc1: q<=8'h20;
	15'h1dc2: q<=8'h22;
	15'h1dc3: q<=8'had;
	15'h1dc4: q<=8'hb8;
	15'h1dc5: q<=8'h50;
	15'h1dc6: q<=8'h06;
	15'h1dc7: q<=8'hca;
	15'h1dc8: q<=8'ha9;
	15'h1dc9: q<=8'h00;
	15'h1dca: q<=8'h9d;
	15'h1dcb: q<=8'h06;
	15'h1dcc: q<=8'h06;
	15'h1dcd: q<=8'h60;
	15'h1dce: q<=8'h48;
	15'h1dcf: q<=8'ha5;
	15'h1dd0: q<=8'h50;
	15'h1dd1: q<=8'h0a;
	15'h1dd2: q<=8'h0a;
	15'h1dd3: q<=8'h0a;
	15'h1dd4: q<=8'h18;
	15'h1dd5: q<=8'h65;
	15'h1dd6: q<=8'h51;
	15'h1dd7: q<=8'h85;
	15'h1dd8: q<=8'h51;
	15'h1dd9: q<=8'h68;
	15'h1dda: q<=8'ha4;
	15'h1ddb: q<=8'h50;
	15'h1ddc: q<=8'h30;
	15'h1ddd: q<=8'h05;
	15'h1dde: q<=8'h69;
	15'h1ddf: q<=8'h00;
	15'h1de0: q<=8'hb8;
	15'h1de1: q<=8'h50;
	15'h1de2: q<=8'h02;
	15'h1de3: q<=8'h69;
	15'h1de4: q<=8'hff;
	15'h1de5: q<=8'ha0;
	15'h1de6: q<=8'h00;
	15'h1de7: q<=8'h84;
	15'h1de8: q<=8'h50;
	15'h1de9: q<=8'h60;
	15'h1dea: q<=8'h20;
	15'h1deb: q<=8'hb4;
	15'h1dec: q<=8'ha8;
	15'h1ded: q<=8'ha9;
	15'h1dee: q<=8'hc0;
	15'h1def: q<=8'ha2;
	15'h1df0: q<=8'h02;
	15'h1df1: q<=8'h20;
	15'h1df2: q<=8'h17;
	15'h1df3: q<=8'hab;
	15'h1df4: q<=8'hce;
	15'h1df5: q<=8'h6e;
	15'h1df6: q<=8'h01;
	15'h1df7: q<=8'h20;
	15'h1df8: q<=8'h97;
	15'h1df9: q<=8'haa;
	15'h1dfa: q<=8'ha2;
	15'h1dfb: q<=8'h0a;
	15'h1dfc: q<=8'h20;
	15'h1dfd: q<=8'h14;
	15'h1dfe: q<=8'hab;
	15'h1dff: q<=8'ha9;
	15'h1e00: q<=8'ha6;
	15'h1e01: q<=8'ha2;
	15'h1e02: q<=8'h0c;
	15'h1e03: q<=8'h20;
	15'h1e04: q<=8'h17;
	15'h1e05: q<=8'hab;
	15'h1e06: q<=8'ha9;
	15'h1e07: q<=8'h9c;
	15'h1e08: q<=8'ha2;
	15'h1e09: q<=8'h0e;
	15'h1e0a: q<=8'h20;
	15'h1e0b: q<=8'h17;
	15'h1e0c: q<=8'hab;
	15'h1e0d: q<=8'ha2;
	15'h1e0e: q<=8'h2c;
	15'h1e0f: q<=8'h20;
	15'h1e10: q<=8'h14;
	15'h1e11: q<=8'hab;
	15'h1e12: q<=8'had;
	15'h1e13: q<=8'h02;
	15'h1e14: q<=8'h06;
	15'h1e15: q<=8'h38;
	15'h1e16: q<=8'hed;
	15'h1e17: q<=8'h04;
	15'h1e18: q<=8'h06;
	15'h1e19: q<=8'h4c;
	15'h1e1a: q<=8'h4e;
	15'h1e1b: q<=8'hae;
	15'h1e1c: q<=8'h20;
	15'h1e1d: q<=8'hb4;
	15'h1e1e: q<=8'ha8;
	15'h1e1f: q<=8'h78;
	15'h1e20: q<=8'had;
	15'h1e21: q<=8'hca;
	15'h1e22: q<=8'h60;
	15'h1e23: q<=8'hac;
	15'h1e24: q<=8'hca;
	15'h1e25: q<=8'h60;
	15'h1e26: q<=8'h84;
	15'h1e27: q<=8'h29;
	15'h1e28: q<=8'h4a;
	15'h1e29: q<=8'h4a;
	15'h1e2a: q<=8'h4a;
	15'h1e2b: q<=8'h4a;
	15'h1e2c: q<=8'h45;
	15'h1e2d: q<=8'h29;
	15'h1e2e: q<=8'h85;
	15'h1e2f: q<=8'h29;
	15'h1e30: q<=8'had;
	15'h1e31: q<=8'hda;
	15'h1e32: q<=8'h60;
	15'h1e33: q<=8'hac;
	15'h1e34: q<=8'hda;
	15'h1e35: q<=8'h60;
	15'h1e36: q<=8'h58;
	15'h1e37: q<=8'h45;
	15'h1e38: q<=8'h29;
	15'h1e39: q<=8'h29;
	15'h1e3a: q<=8'hf0;
	15'h1e3b: q<=8'h45;
	15'h1e3c: q<=8'h29;
	15'h1e3d: q<=8'h85;
	15'h1e3e: q<=8'h29;
	15'h1e3f: q<=8'h98;
	15'h1e40: q<=8'h0a;
	15'h1e41: q<=8'h0a;
	15'h1e42: q<=8'h0a;
	15'h1e43: q<=8'h0a;
	15'h1e44: q<=8'h45;
	15'h1e45: q<=8'h29;
	15'h1e46: q<=8'h8d;
	15'h1e47: q<=8'h1f;
	15'h1e48: q<=8'h01;
	15'h1e49: q<=8'h20;
	15'h1e4a: q<=8'h26;
	15'h1e4b: q<=8'haf;
	15'h1e4c: q<=8'ha9;
	15'h1e4d: q<=8'hff;
	15'h1e4e: q<=8'h85;
	15'h1e4f: q<=8'h63;
	15'h1e50: q<=8'ha2;
	15'h1e51: q<=8'h10;
	15'h1e52: q<=8'h20;
	15'h1e53: q<=8'h14;
	15'h1e54: q<=8'hab;
	15'h1e55: q<=8'ha9;
	15'h1e56: q<=8'h01;
	15'h1e57: q<=8'h85;
	15'h1e58: q<=8'h61;
	15'h1e59: q<=8'h20;
	15'h1e5a: q<=8'hdd;
	15'h1e5b: q<=8'hb0;
	15'h1e5c: q<=8'ha9;
	15'h1e5d: q<=8'h28;
	15'h1e5e: q<=8'h85;
	15'h1e5f: q<=8'h2c;
	15'h1e60: q<=8'ha2;
	15'h1e61: q<=8'h15;
	15'h1e62: q<=8'h86;
	15'h1e63: q<=8'h37;
	15'h1e64: q<=8'h20;
	15'h1e65: q<=8'h0d;
	15'h1e66: q<=8'hab;
	15'h1e67: q<=8'ha9;
	15'h1e68: q<=8'h00;
	15'h1e69: q<=8'h85;
	15'h1e6a: q<=8'h73;
	15'h1e6b: q<=8'ha5;
	15'h1e6c: q<=8'h2c;
	15'h1e6d: q<=8'haa;
	15'h1e6e: q<=8'h38;
	15'h1e6f: q<=8'he9;
	15'h1e70: q<=8'h0a;
	15'h1e71: q<=8'h85;
	15'h1e72: q<=8'h2c;
	15'h1e73: q<=8'ha9;
	15'h1e74: q<=8'hd0;
	15'h1e75: q<=8'h20;
	15'h1e76: q<=8'h75;
	15'h1e77: q<=8'hdf;
	15'h1e78: q<=8'ha0;
	15'h1e79: q<=8'h07;
	15'h1e7a: q<=8'ha5;
	15'h1e7b: q<=8'h63;
	15'h1e7c: q<=8'hc5;
	15'h1e7d: q<=8'h37;
	15'h1e7e: q<=8'hd0;
	15'h1e7f: q<=8'h02;
	15'h1e80: q<=8'ha0;
	15'h1e81: q<=8'h00;
	15'h1e82: q<=8'h20;
	15'h1e83: q<=8'hd1;
	15'h1e84: q<=8'hb0;
	15'h1e85: q<=8'ha9;
	15'h1e86: q<=8'h61;
	15'h1e87: q<=8'ha0;
	15'h1e88: q<=8'h01;
	15'h1e89: q<=8'h20;
	15'h1e8a: q<=8'hb1;
	15'h1e8b: q<=8'hdf;
	15'h1e8c: q<=8'ha9;
	15'h1e8d: q<=8'ha0;
	15'h1e8e: q<=8'h20;
	15'h1e8f: q<=8'h6a;
	15'h1e90: q<=8'hb5;
	15'h1e91: q<=8'ha9;
	15'h1e92: q<=8'h00;
	15'h1e93: q<=8'h85;
	15'h1e94: q<=8'h73;
	15'h1e95: q<=8'haa;
	15'h1e96: q<=8'ha9;
	15'h1e97: q<=8'h08;
	15'h1e98: q<=8'h20;
	15'h1e99: q<=8'h75;
	15'h1e9a: q<=8'hdf;
	15'h1e9b: q<=8'he6;
	15'h1e9c: q<=8'h61;
	15'h1e9d: q<=8'ha5;
	15'h1e9e: q<=8'h37;
	15'h1e9f: q<=8'h20;
	15'h1ea0: q<=8'hf8;
	15'h1ea1: q<=8'hae;
	15'h1ea2: q<=8'ha2;
	15'h1ea3: q<=8'h00;
	15'h1ea4: q<=8'ha9;
	15'h1ea5: q<=8'h08;
	15'h1ea6: q<=8'h20;
	15'h1ea7: q<=8'h75;
	15'h1ea8: q<=8'hdf;
	15'h1ea9: q<=8'ha6;
	15'h1eaa: q<=8'h37;
	15'h1eab: q<=8'hbd;
	15'h1eac: q<=8'h06;
	15'h1ead: q<=8'h07;
	15'h1eae: q<=8'h85;
	15'h1eaf: q<=8'h56;
	15'h1eb0: q<=8'hbd;
	15'h1eb1: q<=8'h07;
	15'h1eb2: q<=8'h07;
	15'h1eb3: q<=8'h85;
	15'h1eb4: q<=8'h57;
	15'h1eb5: q<=8'hbd;
	15'h1eb6: q<=8'h08;
	15'h1eb7: q<=8'h07;
	15'h1eb8: q<=8'h85;
	15'h1eb9: q<=8'h58;
	15'h1eba: q<=8'ha9;
	15'h1ebb: q<=8'h56;
	15'h1ebc: q<=8'ha0;
	15'h1ebd: q<=8'h03;
	15'h1ebe: q<=8'h20;
	15'h1ebf: q<=8'hb1;
	15'h1ec0: q<=8'hdf;
	15'h1ec1: q<=8'hc6;
	15'h1ec2: q<=8'h37;
	15'h1ec3: q<=8'hc6;
	15'h1ec4: q<=8'h37;
	15'h1ec5: q<=8'hc6;
	15'h1ec6: q<=8'h37;
	15'h1ec7: q<=8'h10;
	15'h1ec8: q<=8'h9b;
	15'h1ec9: q<=8'h60;
	15'h1eca: q<=8'had;
	15'h1ecb: q<=8'h56;
	15'h1ecc: q<=8'h01;
	15'h1ecd: q<=8'hf0;
	15'h1ece: q<=8'h14;
	15'h1ecf: q<=8'h85;
	15'h1ed0: q<=8'h58;
	15'h1ed1: q<=8'ha2;
	15'h1ed2: q<=8'h34;
	15'h1ed3: q<=8'h20;
	15'h1ed4: q<=8'h14;
	15'h1ed5: q<=8'hab;
	15'h1ed6: q<=8'ha9;
	15'h1ed7: q<=8'h00;
	15'h1ed8: q<=8'h85;
	15'h1ed9: q<=8'h56;
	15'h1eda: q<=8'h85;
	15'h1edb: q<=8'h57;
	15'h1edc: q<=8'ha9;
	15'h1edd: q<=8'h56;
	15'h1ede: q<=8'ha0;
	15'h1edf: q<=8'h03;
	15'h1ee0: q<=8'h20;
	15'h1ee1: q<=8'hb1;
	15'h1ee2: q<=8'hdf;
	15'h1ee3: q<=8'h18;
	15'h1ee4: q<=8'ha0;
	15'h1ee5: q<=8'h10;
	15'h1ee6: q<=8'ha9;
	15'h1ee7: q<=8'h85;
	15'h1ee8: q<=8'h79;
	15'h1ee9: q<=8'h75;
	15'h1eea: q<=8'hd5;
	15'h1eeb: q<=8'h88;
	15'h1eec: q<=8'h10;
	15'h1eed: q<=8'hfa;
	15'h1eee: q<=8'h85;
	15'h1eef: q<=8'hb5;
	15'h1ef0: q<=8'h60;
	15'h1ef1: q<=8'had;
	15'h1ef2: q<=8'h02;
	15'h1ef3: q<=8'h06;
	15'h1ef4: q<=8'h38;
	15'h1ef5: q<=8'hed;
	15'h1ef6: q<=8'h04;
	15'h1ef7: q<=8'h06;
	15'h1ef8: q<=8'h18;
	15'h1ef9: q<=8'h69;
	15'h1efa: q<=8'h02;
	15'h1efb: q<=8'h85;
	15'h1efc: q<=8'h38;
	15'h1efd: q<=8'ha0;
	15'h1efe: q<=8'h00;
	15'h1eff: q<=8'ha9;
	15'h1f00: q<=8'h02;
	15'h1f01: q<=8'h85;
	15'h1f02: q<=8'h39;
	15'h1f03: q<=8'ha6;
	15'h1f04: q<=8'h38;
	15'h1f05: q<=8'hbd;
	15'h1f06: q<=8'h06;
	15'h1f07: q<=8'h06;
	15'h1f08: q<=8'hc9;
	15'h1f09: q<=8'h1e;
	15'h1f0a: q<=8'h90;
	15'h1f0b: q<=8'h02;
	15'h1f0c: q<=8'ha9;
	15'h1f0d: q<=8'h1a;
	15'h1f0e: q<=8'h0a;
	15'h1f0f: q<=8'haa;
	15'h1f10: q<=8'hbd;
	15'h1f11: q<=8'hfa;
	15'h1f12: q<=8'h31;
	15'h1f13: q<=8'h91;
	15'h1f14: q<=8'h74;
	15'h1f15: q<=8'hc8;
	15'h1f16: q<=8'hbd;
	15'h1f17: q<=8'hfb;
	15'h1f18: q<=8'h31;
	15'h1f19: q<=8'h91;
	15'h1f1a: q<=8'h74;
	15'h1f1b: q<=8'hc8;
	15'h1f1c: q<=8'hc6;
	15'h1f1d: q<=8'h38;
	15'h1f1e: q<=8'hc6;
	15'h1f1f: q<=8'h39;
	15'h1f20: q<=8'h10;
	15'h1f21: q<=8'he1;
	15'h1f22: q<=8'h88;
	15'h1f23: q<=8'h4c;
	15'h1f24: q<=8'h5f;
	15'h1f25: q<=8'hdf;
	15'h1f26: q<=8'had;
	15'h1f27: q<=8'h00;
	15'h1f28: q<=8'h06;
	15'h1f29: q<=8'h0d;
	15'h1f2a: q<=8'h01;
	15'h1f2b: q<=8'h06;
	15'h1f2c: q<=8'hf0;
	15'h1f2d: q<=8'h40;
	15'h1f2e: q<=8'ha2;
	15'h1f2f: q<=8'h12;
	15'h1f30: q<=8'h20;
	15'h1f31: q<=8'h14;
	15'h1f32: q<=8'hab;
	15'h1f33: q<=8'ha9;
	15'h1f34: q<=8'h63;
	15'h1f35: q<=8'h20;
	15'h1f36: q<=8'h71;
	15'h1f37: q<=8'haf;
	15'h1f38: q<=8'ha2;
	15'h1f39: q<=8'h00;
	15'h1f3a: q<=8'h20;
	15'h1f3b: q<=8'h3f;
	15'h1f3c: q<=8'haf;
	15'h1f3d: q<=8'ha2;
	15'h1f3e: q<=8'h01;
	15'h1f3f: q<=8'hbd;
	15'h1f40: q<=8'h00;
	15'h1f41: q<=8'h06;
	15'h1f42: q<=8'hf0;
	15'h1f43: q<=8'h2a;
	15'h1f44: q<=8'h48;
	15'h1f45: q<=8'h86;
	15'h1f46: q<=8'h2e;
	15'h1f47: q<=8'ha0;
	15'h1f48: q<=8'h03;
	15'h1f49: q<=8'h20;
	15'h1f4a: q<=8'hd1;
	15'h1f4b: q<=8'hb0;
	15'h1f4c: q<=8'h20;
	15'h1f4d: q<=8'h0d;
	15'h1f4e: q<=8'hab;
	15'h1f4f: q<=8'ha9;
	15'h1f50: q<=8'hd0;
	15'h1f51: q<=8'ha4;
	15'h1f52: q<=8'h2e;
	15'h1f53: q<=8'hbe;
	15'h1f54: q<=8'h6f;
	15'h1f55: q<=8'haf;
	15'h1f56: q<=8'h20;
	15'h1f57: q<=8'h75;
	15'h1f58: q<=8'hdf;
	15'h1f59: q<=8'h68;
	15'h1f5a: q<=8'h20;
	15'h1f5b: q<=8'h71;
	15'h1f5c: q<=8'haf;
	15'h1f5d: q<=8'ha9;
	15'h1f5e: q<=8'ha0;
	15'h1f5f: q<=8'h20;
	15'h1f60: q<=8'h6a;
	15'h1f61: q<=8'hb5;
	15'h1f62: q<=8'ha9;
	15'h1f63: q<=8'h10;
	15'h1f64: q<=8'ha2;
	15'h1f65: q<=8'h04;
	15'h1f66: q<=8'h20;
	15'h1f67: q<=8'h98;
	15'h1f68: q<=8'hab;
	15'h1f69: q<=8'ha6;
	15'h1f6a: q<=8'h2e;
	15'h1f6b: q<=8'h20;
	15'h1f6c: q<=8'h9e;
	15'h1f6d: q<=8'haa;
	15'h1f6e: q<=8'h60;
	15'h1f6f: q<=8'hc0;
	15'h1f70: q<=8'hb0;
	15'h1f71: q<=8'hc9;
	15'h1f72: q<=8'h63;
	15'h1f73: q<=8'h90;
	15'h1f74: q<=8'h02;
	15'h1f75: q<=8'ha9;
	15'h1f76: q<=8'h63;
	15'h1f77: q<=8'h20;
	15'h1f78: q<=8'hf5;
	15'h1f79: q<=8'haa;
	15'h1f7a: q<=8'ha9;
	15'h1f7b: q<=8'h29;
	15'h1f7c: q<=8'ha0;
	15'h1f7d: q<=8'h01;
	15'h1f7e: q<=8'h4c;
	15'h1f7f: q<=8'hb1;
	15'h1f80: q<=8'hdf;
	15'h1f81: q<=8'h20;
	15'h1f82: q<=8'h48;
	15'h1f83: q<=8'hca;
	15'h1f84: q<=8'hce;
	15'h1f85: q<=8'h6e;
	15'h1f86: q<=8'h01;
	15'h1f87: q<=8'ha0;
	15'h1f88: q<=8'h03;
	15'h1f89: q<=8'h20;
	15'h1f8a: q<=8'hd1;
	15'h1f8b: q<=8'hb0;
	15'h1f8c: q<=8'ha9;
	15'h1f8d: q<=8'h01;
	15'h1f8e: q<=8'h85;
	15'h1f8f: q<=8'h72;
	15'h1f90: q<=8'h20;
	15'h1f91: q<=8'h6a;
	15'h1f92: q<=8'hdf;
	15'h1f93: q<=8'ha2;
	15'h1f94: q<=8'h2c;
	15'h1f95: q<=8'ha9;
	15'h1f96: q<=8'h60;
	15'h1f97: q<=8'h20;
	15'h1f98: q<=8'h17;
	15'h1f99: q<=8'hab;
	15'h1f9a: q<=8'h20;
	15'h1f9b: q<=8'h92;
	15'h1f9c: q<=8'haa;
	15'h1f9d: q<=8'ha2;
	15'h1f9e: q<=8'h07;
	15'h1f9f: q<=8'h86;
	15'h1fa0: q<=8'h37;
	15'h1fa1: q<=8'ha4;
	15'h1fa2: q<=8'h37;
	15'h1fa3: q<=8'hbe;
	15'h1fa4: q<=8'h9b;
	15'h1fa5: q<=8'hb0;
	15'h1fa6: q<=8'h20;
	15'h1fa7: q<=8'h14;
	15'h1fa8: q<=8'hab;
	15'h1fa9: q<=8'hc6;
	15'h1faa: q<=8'h37;
	15'h1fab: q<=8'h10;
	15'h1fac: q<=8'hf4;
	15'h1fad: q<=8'had;
	15'h1fae: q<=8'h00;
	15'h1faf: q<=8'h02;
	15'h1fb0: q<=8'h38;
	15'h1fb1: q<=8'he5;
	15'h1fb2: q<=8'h7b;
	15'h1fb3: q<=8'h10;
	15'h1fb4: q<=8'h07;
	15'h1fb5: q<=8'hc6;
	15'h1fb6: q<=8'h7b;
	15'h1fb7: q<=8'hc6;
	15'h1fb8: q<=8'h7c;
	15'h1fb9: q<=8'hb8;
	15'h1fba: q<=8'h50;
	15'h1fbb: q<=8'h25;
	15'h1fbc: q<=8'hd0;
	15'h1fbd: q<=8'h0d;
	15'h1fbe: q<=8'hc6;
	15'h1fbf: q<=8'h7c;
	15'h1fc0: q<=8'hc6;
	15'h1fc1: q<=8'h7b;
	15'h1fc2: q<=8'h10;
	15'h1fc3: q<=8'h04;
	15'h1fc4: q<=8'he6;
	15'h1fc5: q<=8'h7b;
	15'h1fc6: q<=8'he6;
	15'h1fc7: q<=8'h7c;
	15'h1fc8: q<=8'hb8;
	15'h1fc9: q<=8'h50;
	15'h1fca: q<=8'h16;
	15'h1fcb: q<=8'ha5;
	15'h1fcc: q<=8'h7c;
	15'h1fcd: q<=8'hcd;
	15'h1fce: q<=8'h27;
	15'h1fcf: q<=8'h01;
	15'h1fd0: q<=8'hf0;
	15'h1fd1: q<=8'h02;
	15'h1fd2: q<=8'hb0;
	15'h1fd3: q<=8'h0d;
	15'h1fd4: q<=8'h38;
	15'h1fd5: q<=8'hed;
	15'h1fd6: q<=8'h00;
	15'h1fd7: q<=8'h02;
	15'h1fd8: q<=8'hd0;
	15'h1fd9: q<=8'h01;
	15'h1fda: q<=8'h18;
	15'h1fdb: q<=8'hb0;
	15'h1fdc: q<=8'h04;
	15'h1fdd: q<=8'he6;
	15'h1fde: q<=8'h7b;
	15'h1fdf: q<=8'he6;
	15'h1fe0: q<=8'h7c;
	15'h1fe1: q<=8'ha5;
	15'h1fe2: q<=8'h7c;
	15'h1fe3: q<=8'h85;
	15'h1fe4: q<=8'h3a;
	15'h1fe5: q<=8'ha2;
	15'h1fe6: q<=8'h04;
	15'h1fe7: q<=8'h86;
	15'h1fe8: q<=8'h37;
	15'h1fe9: q<=8'ha0;
	15'h1fea: q<=8'h05;
	15'h1feb: q<=8'h20;
	15'h1fec: q<=8'hd1;
	15'h1fed: q<=8'hb0;
	15'h1fee: q<=8'ha9;
	15'h1fef: q<=8'h00;
	15'h1ff0: q<=8'h85;
	15'h1ff1: q<=8'h73;
	15'h1ff2: q<=8'h20;
	15'h1ff3: q<=8'h0d;
	15'h1ff4: q<=8'hab;
	15'h1ff5: q<=8'ha2;
	15'h1ff6: q<=8'hd8;
	15'h1ff7: q<=8'ha4;
	15'h1ff8: q<=8'h37;
	15'h1ff9: q<=8'hb9;
	15'h1ffa: q<=8'h96;
	15'h1ffb: q<=8'hb0;
	15'h1ffc: q<=8'h18;
	15'h1ffd: q<=8'h69;
	15'h1ffe: q<=8'hf8;
	15'h1fff: q<=8'h20;
	15'h2000: q<=8'h75;
	15'h2001: q<=8'hdf;
	15'h2002: q<=8'ha6;
	15'h2003: q<=8'h3a;
	15'h2004: q<=8'hbc;
	15'h2005: q<=8'hfe;
	15'h2006: q<=8'h91;
	15'h2007: q<=8'hc0;
	15'h2008: q<=8'h63;
	15'h2009: q<=8'hb0;
	15'h200a: q<=8'h37;
	15'h200b: q<=8'hc8;
	15'h200c: q<=8'h98;
	15'h200d: q<=8'h20;
	15'h200e: q<=8'h77;
	15'h200f: q<=8'haf;
	15'h2010: q<=8'ha0;
	15'h2011: q<=8'h03;
	15'h2012: q<=8'h20;
	15'h2013: q<=8'hd1;
	15'h2014: q<=8'hb0;
	15'h2015: q<=8'h20;
	15'h2016: q<=8'h0d;
	15'h2017: q<=8'hab;
	15'h2018: q<=8'ha2;
	15'h2019: q<=8'hba;
	15'h201a: q<=8'ha4;
	15'h201b: q<=8'h37;
	15'h201c: q<=8'hb9;
	15'h201d: q<=8'h96;
	15'h201e: q<=8'hb0;
	15'h201f: q<=8'h18;
	15'h2020: q<=8'h69;
	15'h2021: q<=8'hec;
	15'h2022: q<=8'h20;
	15'h2023: q<=8'h75;
	15'h2024: q<=8'hdf;
	15'h2025: q<=8'ha6;
	15'h2026: q<=8'h3a;
	15'h2027: q<=8'h20;
	15'h2028: q<=8'hc6;
	15'h2029: q<=8'hb0;
	15'h202a: q<=8'h20;
	15'h202b: q<=8'h0d;
	15'h202c: q<=8'hab;
	15'h202d: q<=8'ha2;
	15'h202e: q<=8'hcc;
	15'h202f: q<=8'ha4;
	15'h2030: q<=8'h37;
	15'h2031: q<=8'hb9;
	15'h2032: q<=8'h96;
	15'h2033: q<=8'hb0;
	15'h2034: q<=8'h18;
	15'h2035: q<=8'h69;
	15'h2036: q<=8'h00;
	15'h2037: q<=8'h20;
	15'h2038: q<=8'h75;
	15'h2039: q<=8'hdf;
	15'h203a: q<=8'ha6;
	15'h203b: q<=8'h3a;
	15'h203c: q<=8'hbd;
	15'h203d: q<=8'hfe;
	15'h203e: q<=8'h91;
	15'h203f: q<=8'h20;
	15'h2040: q<=8'he1;
	15'h2041: q<=8'hc4;
	15'h2042: q<=8'hc6;
	15'h2043: q<=8'h3a;
	15'h2044: q<=8'hc6;
	15'h2045: q<=8'h37;
	15'h2046: q<=8'h10;
	15'h2047: q<=8'ha1;
	15'h2048: q<=8'ha9;
	15'h2049: q<=8'h00;
	15'h204a: q<=8'h85;
	15'h204b: q<=8'h73;
	15'h204c: q<=8'h20;
	15'h204d: q<=8'h0d;
	15'h204e: q<=8'hab;
	15'h204f: q<=8'ha2;
	15'h2050: q<=8'h1c;
	15'h2051: q<=8'h20;
	15'h2052: q<=8'h14;
	15'h2053: q<=8'hab;
	15'h2054: q<=8'ha9;
	15'h2055: q<=8'h04;
	15'h2056: q<=8'ha0;
	15'h2057: q<=8'h01;
	15'h2058: q<=8'h20;
	15'h2059: q<=8'hb1;
	15'h205a: q<=8'hdf;
	15'h205b: q<=8'ha0;
	15'h205c: q<=8'h00;
	15'h205d: q<=8'h20;
	15'h205e: q<=8'hd1;
	15'h205f: q<=8'hb0;
	15'h2060: q<=8'h20;
	15'h2061: q<=8'h0d;
	15'h2062: q<=8'hab;
	15'h2063: q<=8'ha2;
	15'h2064: q<=8'hb8;
	15'h2065: q<=8'h20;
	15'h2066: q<=8'hab;
	15'h2067: q<=8'hb0;
	15'h2068: q<=8'h38;
	15'h2069: q<=8'he5;
	15'h206a: q<=8'h7b;
	15'h206b: q<=8'ha8;
	15'h206c: q<=8'hb9;
	15'h206d: q<=8'h96;
	15'h206e: q<=8'hb0;
	15'h206f: q<=8'h38;
	15'h2070: q<=8'he9;
	15'h2071: q<=8'h16;
	15'h2072: q<=8'h20;
	15'h2073: q<=8'h75;
	15'h2074: q<=8'hdf;
	15'h2075: q<=8'ha9;
	15'h2076: q<=8'he0;
	15'h2077: q<=8'h85;
	15'h2078: q<=8'h73;
	15'h2079: q<=8'ha2;
	15'h207a: q<=8'h00;
	15'h207b: q<=8'h86;
	15'h207c: q<=8'h38;
	15'h207d: q<=8'ha0;
	15'h207e: q<=8'h03;
	15'h207f: q<=8'h84;
	15'h2080: q<=8'h37;
	15'h2081: q<=8'ha4;
	15'h2082: q<=8'h38;
	15'h2083: q<=8'hb9;
	15'h2084: q<=8'ha3;
	15'h2085: q<=8'hb0;
	15'h2086: q<=8'haa;
	15'h2087: q<=8'hc8;
	15'h2088: q<=8'hb9;
	15'h2089: q<=8'ha3;
	15'h208a: q<=8'hb0;
	15'h208b: q<=8'hc8;
	15'h208c: q<=8'h84;
	15'h208d: q<=8'h38;
	15'h208e: q<=8'h20;
	15'h208f: q<=8'h75;
	15'h2090: q<=8'hdf;
	15'h2091: q<=8'hc6;
	15'h2092: q<=8'h37;
	15'h2093: q<=8'h10;
	15'h2094: q<=8'hec;
	15'h2095: q<=8'h60;
	15'h2096: q<=8'hbe;
	15'h2097: q<=8'he3;
	15'h2098: q<=8'h09;
	15'h2099: q<=8'h30;
	15'h209a: q<=8'h58;
	15'h209b: q<=8'h14;
	15'h209c: q<=8'h0c;
	15'h209d: q<=8'h0e;
	15'h209e: q<=8'h16;
	15'h209f: q<=8'h18;
	15'h20a0: q<=8'h1e;
	15'h20a1: q<=8'h20;
	15'h20a2: q<=8'h1a;
	15'h20a3: q<=8'h00;
	15'h20a4: q<=8'h26;
	15'h20a5: q<=8'h28;
	15'h20a6: q<=8'h00;
	15'h20a7: q<=8'h00;
	15'h20a8: q<=8'hda;
	15'h20a9: q<=8'hd8;
	15'h20aa: q<=8'h00;
	15'h20ab: q<=8'had;
	15'h20ac: q<=8'h00;
	15'h20ad: q<=8'h02;
	15'h20ae: q<=8'h20;
	15'h20af: q<=8'hce;
	15'h20b0: q<=8'had;
	15'h20b1: q<=8'ha8;
	15'h20b2: q<=8'h10;
	15'h20b3: q<=8'h05;
	15'h20b4: q<=8'ha9;
	15'h20b5: q<=8'h00;
	15'h20b6: q<=8'hb8;
	15'h20b7: q<=8'h50;
	15'h20b8: q<=8'h08;
	15'h20b9: q<=8'hcd;
	15'h20ba: q<=8'h27;
	15'h20bb: q<=8'h01;
	15'h20bc: q<=8'h90;
	15'h20bd: q<=8'h03;
	15'h20be: q<=8'had;
	15'h20bf: q<=8'h27;
	15'h20c0: q<=8'h01;
	15'h20c1: q<=8'h8d;
	15'h20c2: q<=8'h00;
	15'h20c3: q<=8'h02;
	15'h20c4: q<=8'ha8;
	15'h20c5: q<=8'h60;
	15'h20c6: q<=8'h8a;
	15'h20c7: q<=8'h20;
	15'h20c8: q<=8'hb5;
	15'h20c9: q<=8'h91;
	15'h20ca: q<=8'ha9;
	15'h20cb: q<=8'h29;
	15'h20cc: q<=8'ha0;
	15'h20cd: q<=8'h03;
	15'h20ce: q<=8'h4c;
	15'h20cf: q<=8'hb1;
	15'h20d0: q<=8'hdf;
	15'h20d1: q<=8'hc4;
	15'h20d2: q<=8'h9e;
	15'h20d3: q<=8'hf0;
	15'h20d4: q<=8'h07;
	15'h20d5: q<=8'h84;
	15'h20d6: q<=8'h9e;
	15'h20d7: q<=8'ha9;
	15'h20d8: q<=8'h08;
	15'h20d9: q<=8'h4c;
	15'h20da: q<=8'h4c;
	15'h20db: q<=8'hdf;
	15'h20dc: q<=8'h60;
	15'h20dd: q<=8'hc5;
	15'h20de: q<=8'h72;
	15'h20df: q<=8'hf0;
	15'h20e0: q<=8'h05;
	15'h20e1: q<=8'h85;
	15'h20e2: q<=8'h72;
	15'h20e3: q<=8'h4c;
	15'h20e4: q<=8'h6a;
	15'h20e5: q<=8'hdf;
	15'h20e6: q<=8'h60;
	15'h20e7: q<=8'ha9;
	15'h20e8: q<=8'h0a;
	15'h20e9: q<=8'h85;
	15'h20ea: q<=8'h00;
	15'h20eb: q<=8'ha9;
	15'h20ec: q<=8'h00;
	15'h20ed: q<=8'h85;
	15'h20ee: q<=8'h02;
	15'h20ef: q<=8'ha9;
	15'h20f0: q<=8'hdf;
	15'h20f1: q<=8'h85;
	15'h20f2: q<=8'h04;
	15'h20f3: q<=8'ha9;
	15'h20f4: q<=8'h12;
	15'h20f5: q<=8'h85;
	15'h20f6: q<=8'h01;
	15'h20f7: q<=8'ha9;
	15'h20f8: q<=8'h19;
	15'h20f9: q<=8'h8d;
	15'h20fa: q<=8'h4e;
	15'h20fb: q<=8'h01;
	15'h20fc: q<=8'ha9;
	15'h20fd: q<=8'h18;
	15'h20fe: q<=8'h8d;
	15'h20ff: q<=8'h4d;
	15'h2100: q<=8'h01;
	15'h2101: q<=8'h60;
	15'h2102: q<=8'ha9;
	15'h2103: q<=8'h34;
	15'h2104: q<=8'ha2;
	15'h2105: q<=8'haa;
	15'h2106: q<=8'h20;
	15'h2107: q<=8'h5a;
	15'h2108: q<=8'hb1;
	15'h2109: q<=8'had;
	15'h210a: q<=8'h4e;
	15'h210b: q<=8'h01;
	15'h210c: q<=8'hc9;
	15'h210d: q<=8'ha0;
	15'h210e: q<=8'hb0;
	15'h210f: q<=8'h05;
	15'h2110: q<=8'h69;
	15'h2111: q<=8'h14;
	15'h2112: q<=8'h8d;
	15'h2113: q<=8'h4e;
	15'h2114: q<=8'h01;
	15'h2115: q<=8'hc9;
	15'h2116: q<=8'h50;
	15'h2117: q<=8'h90;
	15'h2118: q<=8'h17;
	15'h2119: q<=8'had;
	15'h211a: q<=8'h4d;
	15'h211b: q<=8'h01;
	15'h211c: q<=8'h18;
	15'h211d: q<=8'h69;
	15'h211e: q<=8'h08;
	15'h211f: q<=8'h8d;
	15'h2120: q<=8'h4d;
	15'h2121: q<=8'h01;
	15'h2122: q<=8'hcd;
	15'h2123: q<=8'h4e;
	15'h2124: q<=8'h01;
	15'h2125: q<=8'h90;
	15'h2126: q<=8'h09;
	15'h2127: q<=8'ha9;
	15'h2128: q<=8'ha0;
	15'h2129: q<=8'h8d;
	15'h212a: q<=8'h4d;
	15'h212b: q<=8'h01;
	15'h212c: q<=8'ha9;
	15'h212d: q<=8'h14;
	15'h212e: q<=8'h85;
	15'h212f: q<=8'h01;
	15'h2130: q<=8'h60;
	15'h2131: q<=8'ha9;
	15'h2132: q<=8'h3f;
	15'h2133: q<=8'ha2;
	15'h2134: q<=8'h4e;
	15'h2135: q<=8'h20;
	15'h2136: q<=8'h5a;
	15'h2137: q<=8'hb1;
	15'h2138: q<=8'had;
	15'h2139: q<=8'h4d;
	15'h213a: q<=8'h01;
	15'h213b: q<=8'hc9;
	15'h213c: q<=8'h30;
	15'h213d: q<=8'h90;
	15'h213e: q<=8'h05;
	15'h213f: q<=8'he9;
	15'h2140: q<=8'h01;
	15'h2141: q<=8'h8d;
	15'h2142: q<=8'h4d;
	15'h2143: q<=8'h01;
	15'h2144: q<=8'hc9;
	15'h2145: q<=8'h80;
	15'h2146: q<=8'hb0;
	15'h2147: q<=8'h11;
	15'h2148: q<=8'had;
	15'h2149: q<=8'h4e;
	15'h214a: q<=8'h01;
	15'h214b: q<=8'h38;
	15'h214c: q<=8'he9;
	15'h214d: q<=8'h01;
	15'h214e: q<=8'hcd;
	15'h214f: q<=8'h4d;
	15'h2150: q<=8'h01;
	15'h2151: q<=8'hb0;
	15'h2152: q<=8'h03;
	15'h2153: q<=8'had;
	15'h2154: q<=8'h4d;
	15'h2155: q<=8'h01;
	15'h2156: q<=8'h8d;
	15'h2157: q<=8'h4e;
	15'h2158: q<=8'h01;
	15'h2159: q<=8'h60;
	15'h215a: q<=8'h85;
	15'h215b: q<=8'h57;
	15'h215c: q<=8'h86;
	15'h215d: q<=8'h56;
	15'h215e: q<=8'had;
	15'h215f: q<=8'h4d;
	15'h2160: q<=8'h01;
	15'h2161: q<=8'h85;
	15'h2162: q<=8'h37;
	15'h2163: q<=8'hce;
	15'h2164: q<=8'h6e;
	15'h2165: q<=8'h01;
	15'h2166: q<=8'ha5;
	15'h2167: q<=8'h37;
	15'h2168: q<=8'h0a;
	15'h2169: q<=8'h0a;
	15'h216a: q<=8'h29;
	15'h216b: q<=8'h7f;
	15'h216c: q<=8'ha8;
	15'h216d: q<=8'ha5;
	15'h216e: q<=8'h37;
	15'h216f: q<=8'h4a;
	15'h2170: q<=8'h4a;
	15'h2171: q<=8'h4a;
	15'h2172: q<=8'h4a;
	15'h2173: q<=8'h4a;
	15'h2174: q<=8'h20;
	15'h2175: q<=8'h6c;
	15'h2176: q<=8'hdf;
	15'h2177: q<=8'ha5;
	15'h2178: q<=8'h37;
	15'h2179: q<=8'hcd;
	15'h217a: q<=8'h4d;
	15'h217b: q<=8'h01;
	15'h217c: q<=8'hd0;
	15'h217d: q<=8'h05;
	15'h217e: q<=8'ha9;
	15'h217f: q<=8'h00;
	15'h2180: q<=8'hb8;
	15'h2181: q<=8'h50;
	15'h2182: q<=8'h0c;
	15'h2183: q<=8'h4a;
	15'h2184: q<=8'h4a;
	15'h2185: q<=8'h4a;
	15'h2186: q<=8'hea;
	15'h2187: q<=8'h29;
	15'h2188: q<=8'h07;
	15'h2189: q<=8'hc9;
	15'h218a: q<=8'h07;
	15'h218b: q<=8'hd0;
	15'h218c: q<=8'h02;
	15'h218d: q<=8'ha9;
	15'h218e: q<=8'h03;
	15'h218f: q<=8'ha8;
	15'h2190: q<=8'ha9;
	15'h2191: q<=8'h68;
	15'h2192: q<=8'h20;
	15'h2193: q<=8'h4c;
	15'h2194: q<=8'hdf;
	15'h2195: q<=8'ha5;
	15'h2196: q<=8'h57;
	15'h2197: q<=8'ha6;
	15'h2198: q<=8'h56;
	15'h2199: q<=8'h20;
	15'h219a: q<=8'h39;
	15'h219b: q<=8'hdf;
	15'h219c: q<=8'ha5;
	15'h219d: q<=8'h37;
	15'h219e: q<=8'h18;
	15'h219f: q<=8'h69;
	15'h21a0: q<=8'h02;
	15'h21a1: q<=8'h85;
	15'h21a2: q<=8'h37;
	15'h21a3: q<=8'hcd;
	15'h21a4: q<=8'h4e;
	15'h21a5: q<=8'h01;
	15'h21a6: q<=8'h90;
	15'h21a7: q<=8'hbe;
	15'h21a8: q<=8'ha2;
	15'h21a9: q<=8'h2c;
	15'h21aa: q<=8'ha9;
	15'h21ab: q<=8'hd0;
	15'h21ac: q<=8'h20;
	15'h21ad: q<=8'h17;
	15'h21ae: q<=8'hab;
	15'h21af: q<=8'ha9;
	15'h21b0: q<=8'h3f;
	15'h21b1: q<=8'ha2;
	15'h21b2: q<=8'hf2;
	15'h21b3: q<=8'h4c;
	15'h21b4: q<=8'h39;
	15'h21b5: q<=8'hdf;
	15'h21b6: q<=8'h20;
	15'h21b7: q<=8'hc3;
	15'h21b8: q<=8'hc1;
	15'h21b9: q<=8'had;
	15'h21ba: q<=8'h00;
	15'h21bb: q<=8'h20;
	15'h21bc: q<=8'hcd;
	15'h21bd: q<=8'hc6;
	15'h21be: q<=8'hce;
	15'h21bf: q<=8'hd0;
	15'h21c0: q<=8'h06;
	15'h21c1: q<=8'had;
	15'h21c2: q<=8'h33;
	15'h21c3: q<=8'h01;
	15'h21c4: q<=8'hd0;
	15'h21c5: q<=8'h01;
	15'h21c6: q<=8'h60;
	15'h21c7: q<=8'ha5;
	15'h21c8: q<=8'h01;
	15'h21c9: q<=8'hc9;
	15'h21ca: q<=8'h00;
	15'h21cb: q<=8'hf0;
	15'h21cc: q<=8'h3c;
	15'h21cd: q<=8'ha9;
	15'h21ce: q<=8'h00;
	15'h21cf: q<=8'h20;
	15'h21d0: q<=8'hbe;
	15'h21d1: q<=8'hb2;
	15'h21d2: q<=8'h20;
	15'h21d3: q<=8'h32;
	15'h21d4: q<=8'hb3;
	15'h21d5: q<=8'hb0;
	15'h21d6: q<=8'h1e;
	15'h21d7: q<=8'h20;
	15'h21d8: q<=8'h0d;
	15'h21d9: q<=8'hb2;
	15'h21da: q<=8'had;
	15'h21db: q<=8'h6e;
	15'h21dc: q<=8'h01;
	15'h21dd: q<=8'hf0;
	15'h21de: q<=8'h16;
	15'h21df: q<=8'ha0;
	15'h21e0: q<=8'h27;
	15'h21e1: q<=8'ha9;
	15'h21e2: q<=8'h0e;
	15'h21e3: q<=8'h38;
	15'h21e4: q<=8'hf1;
	15'h21e5: q<=8'hb6;
	15'h21e6: q<=8'h88;
	15'h21e7: q<=8'h10;
	15'h21e8: q<=8'hfb;
	15'h21e9: q<=8'ha8;
	15'h21ea: q<=8'hf0;
	15'h21eb: q<=8'h02;
	15'h21ec: q<=8'h49;
	15'h21ed: q<=8'he5;
	15'h21ee: q<=8'hf0;
	15'h21ef: q<=8'h02;
	15'h21f0: q<=8'h49;
	15'h21f1: q<=8'h29;
	15'h21f2: q<=8'h8d;
	15'h21f3: q<=8'h55;
	15'h21f4: q<=8'h04;
	15'h21f5: q<=8'ha9;
	15'h21f6: q<=8'h00;
	15'h21f7: q<=8'h20;
	15'h21f8: q<=8'hfe;
	15'h21f9: q<=8'hb2;
	15'h21fa: q<=8'had;
	15'h21fb: q<=8'hc4;
	15'h21fc: q<=8'hce;
	15'h21fd: q<=8'h8d;
	15'h21fe: q<=8'h00;
	15'h21ff: q<=8'h20;
	15'h2200: q<=8'had;
	15'h2201: q<=8'hc5;
	15'h2202: q<=8'hce;
	15'h2203: q<=8'h8d;
	15'h2204: q<=8'h01;
	15'h2205: q<=8'h20;
	15'h2206: q<=8'hb8;
	15'h2207: q<=8'h50;
	15'h2208: q<=8'h03;
	15'h2209: q<=8'h4c;
	15'h220a: q<=8'h30;
	15'h220b: q<=8'hb2;
	15'h220c: q<=8'h60;
	15'h220d: q<=8'ha6;
	15'h220e: q<=8'h01;
	15'h220f: q<=8'hbd;
	15'h2210: q<=8'h19;
	15'h2211: q<=8'hb2;
	15'h2212: q<=8'h48;
	15'h2213: q<=8'hbd;
	15'h2214: q<=8'h18;
	15'h2215: q<=8'hb2;
	15'h2216: q<=8'h48;
	15'h2217: q<=8'h60;
	15'h2218: q<=8'h2f;
	15'h2219: q<=8'hb2;
	15'h221a: q<=8'h03;
	15'h221b: q<=8'hd8;
	15'h221c: q<=8'hb9;
	15'h221d: q<=8'hb8;
	15'h221e: q<=8'he9;
	15'h221f: q<=8'had;
	15'h2220: q<=8'h80;
	15'h2221: q<=8'haf;
	15'h2222: q<=8'h1b;
	15'h2223: q<=8'hae;
	15'h2224: q<=8'h61;
	15'h2225: q<=8'haa;
	15'h2226: q<=8'h59;
	15'h2227: q<=8'haa;
	15'h2228: q<=8'h6e;
	15'h2229: q<=8'haa;
	15'h222a: q<=8'h01;
	15'h222b: q<=8'hb1;
	15'h222c: q<=8'h30;
	15'h222d: q<=8'hb1;
	15'h222e: q<=8'h78;
	15'h222f: q<=8'haa;
	15'h2230: q<=8'ha9;
	15'h2231: q<=8'h07;
	15'h2232: q<=8'h20;
	15'h2233: q<=8'hbe;
	15'h2234: q<=8'hb2;
	15'h2235: q<=8'h20;
	15'h2236: q<=8'h86;
	15'h2237: q<=8'hb5;
	15'h2238: q<=8'ha9;
	15'h2239: q<=8'h07;
	15'h223a: q<=8'h20;
	15'h223b: q<=8'hfe;
	15'h223c: q<=8'hb2;
	15'h223d: q<=8'ha9;
	15'h223e: q<=8'h04;
	15'h223f: q<=8'h20;
	15'h2240: q<=8'hbe;
	15'h2241: q<=8'hb2;
	15'h2242: q<=8'h20;
	15'h2243: q<=8'h5b;
	15'h2244: q<=8'hb7;
	15'h2245: q<=8'ha9;
	15'h2246: q<=8'h04;
	15'h2247: q<=8'h20;
	15'h2248: q<=8'hfe;
	15'h2249: q<=8'hb2;
	15'h224a: q<=8'ha9;
	15'h224b: q<=8'h03;
	15'h224c: q<=8'h20;
	15'h224d: q<=8'hbe;
	15'h224e: q<=8'hb2;
	15'h224f: q<=8'h20;
	15'h2250: q<=8'had;
	15'h2251: q<=8'hb5;
	15'h2252: q<=8'ha9;
	15'h2253: q<=8'h03;
	15'h2254: q<=8'h20;
	15'h2255: q<=8'hfe;
	15'h2256: q<=8'hb2;
	15'h2257: q<=8'ha9;
	15'h2258: q<=8'h06;
	15'h2259: q<=8'h20;
	15'h225a: q<=8'hbe;
	15'h225b: q<=8'hb2;
	15'h225c: q<=8'h20;
	15'h225d: q<=8'h9a;
	15'h225e: q<=8'hb7;
	15'h225f: q<=8'ha9;
	15'h2260: q<=8'h06;
	15'h2261: q<=8'h20;
	15'h2262: q<=8'hfe;
	15'h2263: q<=8'hb2;
	15'h2264: q<=8'ha9;
	15'h2265: q<=8'h05;
	15'h2266: q<=8'h20;
	15'h2267: q<=8'hbe;
	15'h2268: q<=8'hb2;
	15'h2269: q<=8'h20;
	15'h226a: q<=8'h98;
	15'h226b: q<=8'hb4;
	15'h226c: q<=8'ha9;
	15'h226d: q<=8'h05;
	15'h226e: q<=8'h20;
	15'h226f: q<=8'hfe;
	15'h2270: q<=8'hb2;
	15'h2271: q<=8'ha9;
	15'h2272: q<=8'h00;
	15'h2273: q<=8'h20;
	15'h2274: q<=8'hbe;
	15'h2275: q<=8'hb2;
	15'h2276: q<=8'h20;
	15'h2277: q<=8'hb4;
	15'h2278: q<=8'ha8;
	15'h2279: q<=8'ha5;
	15'h227a: q<=8'h05;
	15'h227b: q<=8'h30;
	15'h227c: q<=8'h0d;
	15'h227d: q<=8'ha9;
	15'h227e: q<=8'hf2;
	15'h227f: q<=8'h18;
	15'h2280: q<=8'ha0;
	15'h2281: q<=8'h27;
	15'h2282: q<=8'h71;
	15'h2283: q<=8'hb6;
	15'h2284: q<=8'h88;
	15'h2285: q<=8'h10;
	15'h2286: q<=8'hfb;
	15'h2287: q<=8'h8d;
	15'h2288: q<=8'h1b;
	15'h2289: q<=8'h01;
	15'h228a: q<=8'ha9;
	15'h228b: q<=8'h00;
	15'h228c: q<=8'h20;
	15'h228d: q<=8'hfe;
	15'h228e: q<=8'hb2;
	15'h228f: q<=8'h20;
	15'h2290: q<=8'h67;
	15'h2291: q<=8'hb3;
	15'h2292: q<=8'ha9;
	15'h2293: q<=8'h01;
	15'h2294: q<=8'h20;
	15'h2295: q<=8'hbe;
	15'h2296: q<=8'hb2;
	15'h2297: q<=8'h20;
	15'h2298: q<=8'hc2;
	15'h2299: q<=8'hc5;
	15'h229a: q<=8'ha9;
	15'h229b: q<=8'h01;
	15'h229c: q<=8'h20;
	15'h229d: q<=8'hfe;
	15'h229e: q<=8'hb2;
	15'h229f: q<=8'ha9;
	15'h22a0: q<=8'h08;
	15'h22a1: q<=8'h20;
	15'h22a2: q<=8'hbe;
	15'h22a3: q<=8'hb2;
	15'h22a4: q<=8'h20;
	15'h22a5: q<=8'h4d;
	15'h22a6: q<=8'hc5;
	15'h22a7: q<=8'ha9;
	15'h22a8: q<=8'h08;
	15'h22a9: q<=8'h20;
	15'h22aa: q<=8'hfe;
	15'h22ab: q<=8'hb2;
	15'h22ac: q<=8'ha9;
	15'h22ad: q<=8'h00;
	15'h22ae: q<=8'h8d;
	15'h22af: q<=8'h14;
	15'h22b0: q<=8'h01;
	15'h22b1: q<=8'had;
	15'h22b2: q<=8'hc2;
	15'h22b3: q<=8'hce;
	15'h22b4: q<=8'h8d;
	15'h22b5: q<=8'h00;
	15'h22b6: q<=8'h20;
	15'h22b7: q<=8'had;
	15'h22b8: q<=8'hc3;
	15'h22b9: q<=8'hce;
	15'h22ba: q<=8'h8d;
	15'h22bb: q<=8'h01;
	15'h22bc: q<=8'h20;
	15'h22bd: q<=8'h60;
	15'h22be: q<=8'haa;
	15'h22bf: q<=8'h0a;
	15'h22c0: q<=8'ha8;
	15'h22c1: q<=8'hbd;
	15'h22c2: q<=8'h15;
	15'h22c3: q<=8'h04;
	15'h22c4: q<=8'hd0;
	15'h22c5: q<=8'h09;
	15'h22c6: q<=8'hbe;
	15'h22c7: q<=8'h7a;
	15'h22c8: q<=8'hce;
	15'h22c9: q<=8'hb9;
	15'h22ca: q<=8'h7b;
	15'h22cb: q<=8'hce;
	15'h22cc: q<=8'hb8;
	15'h22cd: q<=8'h50;
	15'h22ce: q<=8'h06;
	15'h22cf: q<=8'hbe;
	15'h22d0: q<=8'h68;
	15'h22d1: q<=8'hce;
	15'h22d2: q<=8'hb9;
	15'h22d3: q<=8'h69;
	15'h22d4: q<=8'hce;
	15'h22d5: q<=8'h86;
	15'h22d6: q<=8'h74;
	15'h22d7: q<=8'h85;
	15'h22d8: q<=8'h75;
	15'h22d9: q<=8'ha9;
	15'h22da: q<=8'h00;
	15'h22db: q<=8'h85;
	15'h22dc: q<=8'ha9;
	15'h22dd: q<=8'h60;
	15'h22de: q<=8'haa;
	15'h22df: q<=8'h0a;
	15'h22e0: q<=8'ha8;
	15'h22e1: q<=8'hbd;
	15'h22e2: q<=8'h15;
	15'h22e3: q<=8'h04;
	15'h22e4: q<=8'hd0;
	15'h22e5: q<=8'h09;
	15'h22e6: q<=8'hbe;
	15'h22e7: q<=8'h68;
	15'h22e8: q<=8'hce;
	15'h22e9: q<=8'hb9;
	15'h22ea: q<=8'h69;
	15'h22eb: q<=8'hce;
	15'h22ec: q<=8'hb8;
	15'h22ed: q<=8'h50;
	15'h22ee: q<=8'h06;
	15'h22ef: q<=8'hbe;
	15'h22f0: q<=8'h7a;
	15'h22f1: q<=8'hce;
	15'h22f2: q<=8'hb9;
	15'h22f3: q<=8'h7b;
	15'h22f4: q<=8'hce;
	15'h22f5: q<=8'h86;
	15'h22f6: q<=8'h3b;
	15'h22f7: q<=8'h85;
	15'h22f8: q<=8'h3c;
	15'h22f9: q<=8'ha9;
	15'h22fa: q<=8'h00;
	15'h22fb: q<=8'h85;
	15'h22fc: q<=8'ha9;
	15'h22fd: q<=8'h60;
	15'h22fe: q<=8'h48;
	15'h22ff: q<=8'h20;
	15'h2300: q<=8'h09;
	15'h2301: q<=8'hdf;
	15'h2302: q<=8'h68;
	15'h2303: q<=8'haa;
	15'h2304: q<=8'h0a;
	15'h2305: q<=8'ha8;
	15'h2306: q<=8'hb9;
	15'h2307: q<=8'h8c;
	15'h2308: q<=8'hce;
	15'h2309: q<=8'h85;
	15'h230a: q<=8'h3b;
	15'h230b: q<=8'hb9;
	15'h230c: q<=8'h8d;
	15'h230d: q<=8'hce;
	15'h230e: q<=8'h85;
	15'h230f: q<=8'h3c;
	15'h2310: q<=8'hbd;
	15'h2311: q<=8'h15;
	15'h2312: q<=8'h04;
	15'h2313: q<=8'h49;
	15'h2314: q<=8'h01;
	15'h2315: q<=8'h9d;
	15'h2316: q<=8'h15;
	15'h2317: q<=8'h04;
	15'h2318: q<=8'hd0;
	15'h2319: q<=8'h09;
	15'h231a: q<=8'hb9;
	15'h231b: q<=8'h9e;
	15'h231c: q<=8'hce;
	15'h231d: q<=8'hbe;
	15'h231e: q<=8'h9f;
	15'h231f: q<=8'hce;
	15'h2320: q<=8'hb8;
	15'h2321: q<=8'h50;
	15'h2322: q<=8'h06;
	15'h2323: q<=8'hb9;
	15'h2324: q<=8'hb0;
	15'h2325: q<=8'hce;
	15'h2326: q<=8'hbe;
	15'h2327: q<=8'hb1;
	15'h2328: q<=8'hce;
	15'h2329: q<=8'ha0;
	15'h232a: q<=8'h00;
	15'h232b: q<=8'h91;
	15'h232c: q<=8'h3b;
	15'h232d: q<=8'h8a;
	15'h232e: q<=8'hc8;
	15'h232f: q<=8'h91;
	15'h2330: q<=8'h3b;
	15'h2331: q<=8'h60;
	15'h2332: q<=8'had;
	15'h2333: q<=8'hc4;
	15'h2334: q<=8'hce;
	15'h2335: q<=8'hcd;
	15'h2336: q<=8'h00;
	15'h2337: q<=8'h20;
	15'h2338: q<=8'hf0;
	15'h2339: q<=8'h05;
	15'h233a: q<=8'h8d;
	15'h233b: q<=8'h00;
	15'h233c: q<=8'h20;
	15'h233d: q<=8'h38;
	15'h233e: q<=8'h60;
	15'h233f: q<=8'had;
	15'h2340: q<=8'h15;
	15'h2341: q<=8'h04;
	15'h2342: q<=8'hd0;
	15'h2343: q<=8'h05;
	15'h2344: q<=8'ha2;
	15'h2345: q<=8'h02;
	15'h2346: q<=8'hb8;
	15'h2347: q<=8'h50;
	15'h2348: q<=8'h02;
	15'h2349: q<=8'ha2;
	15'h234a: q<=8'h08;
	15'h234b: q<=8'hbd;
	15'h234c: q<=8'h9e;
	15'h234d: q<=8'hce;
	15'h234e: q<=8'ha0;
	15'h234f: q<=8'h00;
	15'h2350: q<=8'h8c;
	15'h2351: q<=8'h6e;
	15'h2352: q<=8'h01;
	15'h2353: q<=8'h91;
	15'h2354: q<=8'h74;
	15'h2355: q<=8'hc8;
	15'h2356: q<=8'hbd;
	15'h2357: q<=8'h9f;
	15'h2358: q<=8'hce;
	15'h2359: q<=8'h91;
	15'h235a: q<=8'h74;
	15'h235b: q<=8'hbd;
	15'h235c: q<=8'h68;
	15'h235d: q<=8'hce;
	15'h235e: q<=8'h85;
	15'h235f: q<=8'h74;
	15'h2360: q<=8'hbd;
	15'h2361: q<=8'h69;
	15'h2362: q<=8'hce;
	15'h2363: q<=8'h85;
	15'h2364: q<=8'h75;
	15'h2365: q<=8'h18;
	15'h2366: q<=8'h60;
	15'h2367: q<=8'had;
	15'h2368: q<=8'h14;
	15'h2369: q<=8'h01;
	15'h236a: q<=8'hf0;
	15'h236b: q<=8'h0d;
	15'h236c: q<=8'ha9;
	15'h236d: q<=8'h02;
	15'h236e: q<=8'h20;
	15'h236f: q<=8'hbe;
	15'h2370: q<=8'hb2;
	15'h2371: q<=8'h20;
	15'h2372: q<=8'h0d;
	15'h2373: q<=8'hc3;
	15'h2374: q<=8'ha9;
	15'h2375: q<=8'h02;
	15'h2376: q<=8'h20;
	15'h2377: q<=8'hfe;
	15'h2378: q<=8'hb2;
	15'h2379: q<=8'ha9;
	15'h237a: q<=8'h02;
	15'h237b: q<=8'h20;
	15'h237c: q<=8'hde;
	15'h237d: q<=8'hb2;
	15'h237e: q<=8'ha9;
	15'h237f: q<=8'h00;
	15'h2380: q<=8'ha2;
	15'h2381: q<=8'h0f;
	15'h2382: q<=8'h9d;
	15'h2383: q<=8'h25;
	15'h2384: q<=8'h04;
	15'h2385: q<=8'hca;
	15'h2386: q<=8'h10;
	15'h2387: q<=8'hfa;
	15'h2388: q<=8'had;
	15'h2389: q<=8'h06;
	15'h238a: q<=8'h01;
	15'h238b: q<=8'h30;
	15'h238c: q<=8'h49;
	15'h238d: q<=8'hae;
	15'h238e: q<=8'h1c;
	15'h238f: q<=8'h01;
	15'h2390: q<=8'hbd;
	15'h2391: q<=8'hdf;
	15'h2392: q<=8'h02;
	15'h2393: q<=8'hf0;
	15'h2394: q<=8'h3e;
	15'h2395: q<=8'ha0;
	15'h2396: q<=8'h00;
	15'h2397: q<=8'hbd;
	15'h2398: q<=8'h83;
	15'h2399: q<=8'h02;
	15'h239a: q<=8'h29;
	15'h239b: q<=8'h07;
	15'h239c: q<=8'hc9;
	15'h239d: q<=8'h01;
	15'h239e: q<=8'hd0;
	15'h239f: q<=8'h33;
	15'h23a0: q<=8'hc8;
	15'h23a1: q<=8'h84;
	15'h23a2: q<=8'h29;
	15'h23a3: q<=8'hbd;
	15'h23a4: q<=8'h83;
	15'h23a5: q<=8'h02;
	15'h23a6: q<=8'h29;
	15'h23a7: q<=8'h80;
	15'h23a8: q<=8'hd0;
	15'h23a9: q<=8'h1c;
	15'h23aa: q<=8'had;
	15'h23ab: q<=8'h48;
	15'h23ac: q<=8'h01;
	15'h23ad: q<=8'h30;
	15'h23ae: q<=8'h0c;
	15'h23af: q<=8'hbd;
	15'h23b0: q<=8'hdf;
	15'h23b1: q<=8'h02;
	15'h23b2: q<=8'hcd;
	15'h23b3: q<=8'h57;
	15'h23b4: q<=8'h01;
	15'h23b5: q<=8'hb0;
	15'h23b6: q<=8'h04;
	15'h23b7: q<=8'he6;
	15'h23b8: q<=8'h29;
	15'h23b9: q<=8'he6;
	15'h23ba: q<=8'h29;
	15'h23bb: q<=8'ha5;
	15'h23bc: q<=8'h29;
	15'h23bd: q<=8'hbc;
	15'h23be: q<=8'hcc;
	15'h23bf: q<=8'h02;
	15'h23c0: q<=8'h19;
	15'h23c1: q<=8'h25;
	15'h23c2: q<=8'h04;
	15'h23c3: q<=8'h99;
	15'h23c4: q<=8'h25;
	15'h23c5: q<=8'h04;
	15'h23c6: q<=8'hbc;
	15'h23c7: q<=8'hb9;
	15'h23c8: q<=8'h02;
	15'h23c9: q<=8'ha5;
	15'h23ca: q<=8'h29;
	15'h23cb: q<=8'h09;
	15'h23cc: q<=8'h80;
	15'h23cd: q<=8'h19;
	15'h23ce: q<=8'h25;
	15'h23cf: q<=8'h04;
	15'h23d0: q<=8'h99;
	15'h23d1: q<=8'h25;
	15'h23d2: q<=8'h04;
	15'h23d3: q<=8'hca;
	15'h23d4: q<=8'h10;
	15'h23d5: q<=8'hba;
	15'h23d6: q<=8'ha9;
	15'h23d7: q<=8'h06;
	15'h23d8: q<=8'hac;
	15'h23d9: q<=8'h25;
	15'h23da: q<=8'h01;
	15'h23db: q<=8'hf0;
	15'h23dc: q<=8'h0c;
	15'h23dd: q<=8'h30;
	15'h23de: q<=8'h0a;
	15'h23df: q<=8'ha5;
	15'h23e0: q<=8'h03;
	15'h23e1: q<=8'h29;
	15'h23e2: q<=8'h07;
	15'h23e3: q<=8'hc9;
	15'h23e4: q<=8'h07;
	15'h23e5: q<=8'hd0;
	15'h23e6: q<=8'h02;
	15'h23e7: q<=8'ha9;
	15'h23e8: q<=8'h01;
	15'h23e9: q<=8'h85;
	15'h23ea: q<=8'h29;
	15'h23eb: q<=8'ha0;
	15'h23ec: q<=8'hff;
	15'h23ed: q<=8'ha2;
	15'h23ee: q<=8'hff;
	15'h23ef: q<=8'h86;
	15'h23f0: q<=8'h2c;
	15'h23f1: q<=8'had;
	15'h23f2: q<=8'h02;
	15'h23f3: q<=8'h02;
	15'h23f4: q<=8'hf0;
	15'h23f5: q<=8'h0b;
	15'h23f6: q<=8'had;
	15'h23f7: q<=8'h01;
	15'h23f8: q<=8'h02;
	15'h23f9: q<=8'h30;
	15'h23fa: q<=8'h06;
	15'h23fb: q<=8'hae;
	15'h23fc: q<=8'h00;
	15'h23fd: q<=8'h02;
	15'h23fe: q<=8'hac;
	15'h23ff: q<=8'h01;
	15'h2400: q<=8'h02;
	15'h2401: q<=8'h86;
	15'h2402: q<=8'h2a;
	15'h2403: q<=8'h84;
	15'h2404: q<=8'h2b;
	15'h2405: q<=8'had;
	15'h2406: q<=8'h24;
	15'h2407: q<=8'h01;
	15'h2408: q<=8'h30;
	15'h2409: q<=8'h08;
	15'h240a: q<=8'h29;
	15'h240b: q<=8'h0e;
	15'h240c: q<=8'h4a;
	15'h240d: q<=8'h85;
	15'h240e: q<=8'h2c;
	15'h240f: q<=8'hce;
	15'h2410: q<=8'h24;
	15'h2411: q<=8'h01;
	15'h2412: q<=8'ha2;
	15'h2413: q<=8'h0f;
	15'h2414: q<=8'ha0;
	15'h2415: q<=8'h06;
	15'h2416: q<=8'hbd;
	15'h2417: q<=8'h25;
	15'h2418: q<=8'h04;
	15'h2419: q<=8'hf0;
	15'h241a: q<=8'h0c;
	15'h241b: q<=8'h29;
	15'h241c: q<=8'h02;
	15'h241d: q<=8'hf0;
	15'h241e: q<=8'h05;
	15'h241f: q<=8'ha5;
	15'h2420: q<=8'h03;
	15'h2421: q<=8'h29;
	15'h2422: q<=8'h01;
	15'h2423: q<=8'ha8;
	15'h2424: q<=8'hb8;
	15'h2425: q<=8'h50;
	15'h2426: q<=8'h24;
	15'h2427: q<=8'he4;
	15'h2428: q<=8'h2a;
	15'h2429: q<=8'hf0;
	15'h242a: q<=8'h02;
	15'h242b: q<=8'he4;
	15'h242c: q<=8'h2b;
	15'h242d: q<=8'hd0;
	15'h242e: q<=8'h05;
	15'h242f: q<=8'ha0;
	15'h2430: q<=8'h01;
	15'h2431: q<=8'hb8;
	15'h2432: q<=8'h50;
	15'h2433: q<=8'h17;
	15'h2434: q<=8'had;
	15'h2435: q<=8'h24;
	15'h2436: q<=8'h01;
	15'h2437: q<=8'h30;
	15'h2438: q<=8'h10;
	15'h2439: q<=8'h8a;
	15'h243a: q<=8'h18;
	15'h243b: q<=8'h65;
	15'h243c: q<=8'h2c;
	15'h243d: q<=8'h29;
	15'h243e: q<=8'h07;
	15'h243f: q<=8'hc9;
	15'h2440: q<=8'h07;
	15'h2441: q<=8'hd0;
	15'h2442: q<=8'h02;
	15'h2443: q<=8'ha9;
	15'h2444: q<=8'h03;
	15'h2445: q<=8'ha8;
	15'h2446: q<=8'hb8;
	15'h2447: q<=8'h50;
	15'h2448: q<=8'h02;
	15'h2449: q<=8'ha4;
	15'h244a: q<=8'h29;
	15'h244b: q<=8'h98;
	15'h244c: q<=8'hbc;
	15'h244d: q<=8'h76;
	15'h244e: q<=8'hb4;
	15'h244f: q<=8'h91;
	15'h2450: q<=8'h3b;
	15'h2451: q<=8'hca;
	15'h2452: q<=8'h10;
	15'h2453: q<=8'hc0;
	15'h2454: q<=8'ha2;
	15'h2455: q<=8'h0f;
	15'h2456: q<=8'h2c;
	15'h2457: q<=8'h11;
	15'h2458: q<=8'h01;
	15'h2459: q<=8'h10;
	15'h245a: q<=8'h01;
	15'h245b: q<=8'hca;
	15'h245c: q<=8'ha0;
	15'h245d: q<=8'hc0;
	15'h245e: q<=8'hbd;
	15'h245f: q<=8'h25;
	15'h2460: q<=8'h04;
	15'h2461: q<=8'h10;
	15'h2462: q<=8'h02;
	15'h2463: q<=8'ha0;
	15'h2464: q<=8'h00;
	15'h2465: q<=8'h84;
	15'h2466: q<=8'h58;
	15'h2467: q<=8'hbc;
	15'h2468: q<=8'h87;
	15'h2469: q<=8'hb4;
	15'h246a: q<=8'hb1;
	15'h246b: q<=8'hb0;
	15'h246c: q<=8'h29;
	15'h246d: q<=8'h1f;
	15'h246e: q<=8'h05;
	15'h246f: q<=8'h58;
	15'h2470: q<=8'h91;
	15'h2471: q<=8'hb0;
	15'h2472: q<=8'hca;
	15'h2473: q<=8'h10;
	15'h2474: q<=8'he7;
	15'h2475: q<=8'h60;
	15'h2476: q<=8'ha8;
	15'h2477: q<=8'h9c;
	15'h2478: q<=8'h92;
	15'h2479: q<=8'h86;
	15'h247a: q<=8'h7c;
	15'h247b: q<=8'h70;
	15'h247c: q<=8'h66;
	15'h247d: q<=8'h5a;
	15'h247e: q<=8'h50;
	15'h247f: q<=8'h44;
	15'h2480: q<=8'h3a;
	15'h2481: q<=8'h2e;
	15'h2482: q<=8'h24;
	15'h2483: q<=8'h18;
	15'h2484: q<=8'h0e;
	15'h2485: q<=8'h02;
	15'h2486: q<=8'hb2;
	15'h2487: q<=8'h3b;
	15'h2488: q<=8'h37;
	15'h2489: q<=8'h33;
	15'h248a: q<=8'h2f;
	15'h248b: q<=8'h2b;
	15'h248c: q<=8'h27;
	15'h248d: q<=8'h23;
	15'h248e: q<=8'h1f;
	15'h248f: q<=8'h1b;
	15'h2490: q<=8'h17;
	15'h2491: q<=8'h13;
	15'h2492: q<=8'h0f;
	15'h2493: q<=8'h0b;
	15'h2494: q<=8'h07;
	15'h2495: q<=8'h03;
	15'h2496: q<=8'h3f;
	15'h2497: q<=8'h1d;
	15'h2498: q<=8'ha0;
	15'h2499: q<=8'h0c;
	15'h249a: q<=8'h84;
	15'h249b: q<=8'h9e;
	15'h249c: q<=8'ha9;
	15'h249d: q<=8'h08;
	15'h249e: q<=8'h20;
	15'h249f: q<=8'h4c;
	15'h24a0: q<=8'hdf;
	15'h24a1: q<=8'ha2;
	15'h24a2: q<=8'h66;
	15'h24a3: q<=8'h20;
	15'h24a4: q<=8'h65;
	15'h24a5: q<=8'hc7;
	15'h24a6: q<=8'ha9;
	15'h24a7: q<=8'h12;
	15'h24a8: q<=8'h85;
	15'h24a9: q<=8'h56;
	15'h24aa: q<=8'ha2;
	15'h24ab: q<=8'h3f;
	15'h24ac: q<=8'h86;
	15'h24ad: q<=8'h37;
	15'h24ae: q<=8'ha0;
	15'h24af: q<=8'h00;
	15'h24b0: q<=8'ha6;
	15'h24b1: q<=8'h37;
	15'h24b2: q<=8'hbd;
	15'h24b3: q<=8'h43;
	15'h24b4: q<=8'h02;
	15'h24b5: q<=8'hd0;
	15'h24b6: q<=8'h03;
	15'h24b7: q<=8'h4c;
	15'h24b8: q<=8'h49;
	15'h24b9: q<=8'hb5;
	15'h24ba: q<=8'hc9;
	15'h24bb: q<=8'h50;
	15'h24bc: q<=8'h90;
	15'h24bd: q<=8'h02;
	15'h24be: q<=8'hc6;
	15'h24bf: q<=8'h37;
	15'h24c0: q<=8'h48;
	15'h24c1: q<=8'h29;
	15'h24c2: q<=8'h3f;
	15'h24c3: q<=8'h91;
	15'h24c4: q<=8'h74;
	15'h24c5: q<=8'h68;
	15'h24c6: q<=8'h2a;
	15'h24c7: q<=8'h2a;
	15'h24c8: q<=8'h2a;
	15'h24c9: q<=8'h29;
	15'h24ca: q<=8'h03;
	15'h24cb: q<=8'h18;
	15'h24cc: q<=8'h69;
	15'h24cd: q<=8'h01;
	15'h24ce: q<=8'h09;
	15'h24cf: q<=8'h70;
	15'h24d0: q<=8'hc8;
	15'h24d1: q<=8'h91;
	15'h24d2: q<=8'h74;
	15'h24d3: q<=8'hc8;
	15'h24d4: q<=8'hbd;
	15'h24d5: q<=8'h03;
	15'h24d6: q<=8'h02;
	15'h24d7: q<=8'haa;
	15'h24d8: q<=8'hbd;
	15'h24d9: q<=8'h8a;
	15'h24da: q<=8'h03;
	15'h24db: q<=8'h38;
	15'h24dc: q<=8'he5;
	15'h24dd: q<=8'h68;
	15'h24de: q<=8'h85;
	15'h24df: q<=8'h63;
	15'h24e0: q<=8'h91;
	15'h24e1: q<=8'h74;
	15'h24e2: q<=8'hc8;
	15'h24e3: q<=8'hbd;
	15'h24e4: q<=8'h7a;
	15'h24e5: q<=8'h03;
	15'h24e6: q<=8'he5;
	15'h24e7: q<=8'h69;
	15'h24e8: q<=8'h85;
	15'h24e9: q<=8'h64;
	15'h24ea: q<=8'h29;
	15'h24eb: q<=8'h1f;
	15'h24ec: q<=8'h91;
	15'h24ed: q<=8'h74;
	15'h24ee: q<=8'hc8;
	15'h24ef: q<=8'hbd;
	15'h24f0: q<=8'h6a;
	15'h24f1: q<=8'h03;
	15'h24f2: q<=8'h85;
	15'h24f3: q<=8'h61;
	15'h24f4: q<=8'h91;
	15'h24f5: q<=8'h74;
	15'h24f6: q<=8'hc8;
	15'h24f7: q<=8'hbd;
	15'h24f8: q<=8'h5a;
	15'h24f9: q<=8'h03;
	15'h24fa: q<=8'h85;
	15'h24fb: q<=8'h62;
	15'h24fc: q<=8'h29;
	15'h24fd: q<=8'h1f;
	15'h24fe: q<=8'h91;
	15'h24ff: q<=8'h74;
	15'h2500: q<=8'hc8;
	15'h2501: q<=8'ha9;
	15'h2502: q<=8'h00;
	15'h2503: q<=8'h91;
	15'h2504: q<=8'h74;
	15'h2505: q<=8'hc8;
	15'h2506: q<=8'h91;
	15'h2507: q<=8'h74;
	15'h2508: q<=8'hc8;
	15'h2509: q<=8'h91;
	15'h250a: q<=8'h74;
	15'h250b: q<=8'ha9;
	15'h250c: q<=8'ha0;
	15'h250d: q<=8'hc8;
	15'h250e: q<=8'h91;
	15'h250f: q<=8'h74;
	15'h2510: q<=8'hc8;
	15'h2511: q<=8'ha5;
	15'h2512: q<=8'h63;
	15'h2513: q<=8'h49;
	15'h2514: q<=8'hff;
	15'h2515: q<=8'h18;
	15'h2516: q<=8'h69;
	15'h2517: q<=8'h01;
	15'h2518: q<=8'h91;
	15'h2519: q<=8'h74;
	15'h251a: q<=8'hc8;
	15'h251b: q<=8'ha5;
	15'h251c: q<=8'h64;
	15'h251d: q<=8'h49;
	15'h251e: q<=8'hff;
	15'h251f: q<=8'h69;
	15'h2520: q<=8'h00;
	15'h2521: q<=8'h29;
	15'h2522: q<=8'h1f;
	15'h2523: q<=8'h91;
	15'h2524: q<=8'h74;
	15'h2525: q<=8'hc8;
	15'h2526: q<=8'ha5;
	15'h2527: q<=8'h61;
	15'h2528: q<=8'h49;
	15'h2529: q<=8'hff;
	15'h252a: q<=8'h18;
	15'h252b: q<=8'h69;
	15'h252c: q<=8'h01;
	15'h252d: q<=8'h91;
	15'h252e: q<=8'h74;
	15'h252f: q<=8'hc8;
	15'h2530: q<=8'ha5;
	15'h2531: q<=8'h62;
	15'h2532: q<=8'h49;
	15'h2533: q<=8'hff;
	15'h2534: q<=8'h69;
	15'h2535: q<=8'h00;
	15'h2536: q<=8'h29;
	15'h2537: q<=8'h1f;
	15'h2538: q<=8'h91;
	15'h2539: q<=8'h74;
	15'h253a: q<=8'hc8;
	15'h253b: q<=8'hc0;
	15'h253c: q<=8'hf0;
	15'h253d: q<=8'h90;
	15'h253e: q<=8'h06;
	15'h253f: q<=8'h88;
	15'h2540: q<=8'h20;
	15'h2541: q<=8'h5f;
	15'h2542: q<=8'hdf;
	15'h2543: q<=8'ha0;
	15'h2544: q<=8'h00;
	15'h2545: q<=8'hc6;
	15'h2546: q<=8'h56;
	15'h2547: q<=8'h30;
	15'h2548: q<=8'h07;
	15'h2549: q<=8'hc6;
	15'h254a: q<=8'h37;
	15'h254b: q<=8'h30;
	15'h254c: q<=8'h03;
	15'h254d: q<=8'h4c;
	15'h254e: q<=8'hb0;
	15'h254f: q<=8'hb4;
	15'h2550: q<=8'h98;
	15'h2551: q<=8'hf0;
	15'h2552: q<=8'h04;
	15'h2553: q<=8'h88;
	15'h2554: q<=8'h20;
	15'h2555: q<=8'h5f;
	15'h2556: q<=8'hdf;
	15'h2557: q<=8'ha5;
	15'h2558: q<=8'hb5;
	15'h2559: q<=8'hf0;
	15'h255a: q<=8'h0a;
	15'h255b: q<=8'ha5;
	15'h255c: q<=8'h46;
	15'h255d: q<=8'hc9;
	15'h255e: q<=8'h0a;
	15'h255f: q<=8'h90;
	15'h2560: q<=8'h04;
	15'h2561: q<=8'ha9;
	15'h2562: q<=8'h7a;
	15'h2563: q<=8'h85;
	15'h2564: q<=8'h53;
	15'h2565: q<=8'ha9;
	15'h2566: q<=8'h01;
	15'h2567: q<=8'h4c;
	15'h2568: q<=8'h6a;
	15'h2569: q<=8'hdf;
	15'h256a: q<=8'h48;
	15'h256b: q<=8'ha0;
	15'h256c: q<=8'h00;
	15'h256d: q<=8'h98;
	15'h256e: q<=8'h91;
	15'h256f: q<=8'h74;
	15'h2570: q<=8'hc8;
	15'h2571: q<=8'h91;
	15'h2572: q<=8'h74;
	15'h2573: q<=8'hc8;
	15'h2574: q<=8'h91;
	15'h2575: q<=8'h74;
	15'h2576: q<=8'hc8;
	15'h2577: q<=8'h68;
	15'h2578: q<=8'h91;
	15'h2579: q<=8'h74;
	15'h257a: q<=8'ha9;
	15'h257b: q<=8'h04;
	15'h257c: q<=8'h18;
	15'h257d: q<=8'h65;
	15'h257e: q<=8'h74;
	15'h257f: q<=8'h85;
	15'h2580: q<=8'h74;
	15'h2581: q<=8'h90;
	15'h2582: q<=8'h02;
	15'h2583: q<=8'he6;
	15'h2584: q<=8'h75;
	15'h2585: q<=8'h60;
	15'h2586: q<=8'ha9;
	15'h2587: q<=8'h01;
	15'h2588: q<=8'h85;
	15'h2589: q<=8'h9e;
	15'h258a: q<=8'had;
	15'h258b: q<=8'h02;
	15'h258c: q<=8'h02;
	15'h258d: q<=8'hf0;
	15'h258e: q<=8'h1d;
	15'h258f: q<=8'hc9;
	15'h2590: q<=8'hf0;
	15'h2591: q<=8'hb0;
	15'h2592: q<=8'h19;
	15'h2593: q<=8'h85;
	15'h2594: q<=8'h57;
	15'h2595: q<=8'h85;
	15'h2596: q<=8'h2f;
	15'h2597: q<=8'had;
	15'h2598: q<=8'h01;
	15'h2599: q<=8'h02;
	15'h259a: q<=8'hc9;
	15'h259b: q<=8'h81;
	15'h259c: q<=8'hf0;
	15'h259d: q<=8'h0e;
	15'h259e: q<=8'hac;
	15'h259f: q<=8'h00;
	15'h25a0: q<=8'h02;
	15'h25a1: q<=8'ha5;
	15'h25a2: q<=8'h51;
	15'h25a3: q<=8'h4a;
	15'h25a4: q<=8'h29;
	15'h25a5: q<=8'h07;
	15'h25a6: q<=8'h18;
	15'h25a7: q<=8'h69;
	15'h25a8: q<=8'h01;
	15'h25a9: q<=8'h20;
	15'h25aa: q<=8'ha0;
	15'h25ab: q<=8'hbd;
	15'h25ac: q<=8'h60;
	15'h25ad: q<=8'had;
	15'h25ae: q<=8'h06;
	15'h25af: q<=8'h01;
	15'h25b0: q<=8'h30;
	15'h25b1: q<=8'h24;
	15'h25b2: q<=8'ha2;
	15'h25b3: q<=8'h06;
	15'h25b4: q<=8'h86;
	15'h25b5: q<=8'h37;
	15'h25b6: q<=8'ha6;
	15'h25b7: q<=8'h37;
	15'h25b8: q<=8'hbd;
	15'h25b9: q<=8'hdf;
	15'h25ba: q<=8'h02;
	15'h25bb: q<=8'hf0;
	15'h25bc: q<=8'h15;
	15'h25bd: q<=8'h85;
	15'h25be: q<=8'h57;
	15'h25bf: q<=8'hbd;
	15'h25c0: q<=8'h83;
	15'h25c1: q<=8'h02;
	15'h25c2: q<=8'h29;
	15'h25c3: q<=8'h18;
	15'h25c4: q<=8'h4a;
	15'h25c5: q<=8'h4a;
	15'h25c6: q<=8'h4a;
	15'h25c7: q<=8'h85;
	15'h25c8: q<=8'h55;
	15'h25c9: q<=8'hbd;
	15'h25ca: q<=8'h83;
	15'h25cb: q<=8'h02;
	15'h25cc: q<=8'h29;
	15'h25cd: q<=8'h07;
	15'h25ce: q<=8'h0a;
	15'h25cf: q<=8'h20;
	15'h25d0: q<=8'hd7;
	15'h25d1: q<=8'hb5;
	15'h25d2: q<=8'hc6;
	15'h25d3: q<=8'h37;
	15'h25d4: q<=8'h10;
	15'h25d5: q<=8'he0;
	15'h25d6: q<=8'h60;
	15'h25d7: q<=8'ha8;
	15'h25d8: q<=8'hb9;
	15'h25d9: q<=8'he2;
	15'h25da: q<=8'hb5;
	15'h25db: q<=8'h48;
	15'h25dc: q<=8'hb9;
	15'h25dd: q<=8'he1;
	15'h25de: q<=8'hb5;
	15'h25df: q<=8'h48;
	15'h25e0: q<=8'h60;
	15'h25e1: q<=8'hea;
	15'h25e2: q<=8'hb5;
	15'h25e3: q<=8'h1a;
	15'h25e4: q<=8'hb7;
	15'h25e5: q<=8'h0e;
	15'h25e6: q<=8'hb6;
	15'h25e7: q<=8'h21;
	15'h25e8: q<=8'hb6;
	15'h25e9: q<=8'h9a;
	15'h25ea: q<=8'hb6;
	15'h25eb: q<=8'ha9;
	15'h25ec: q<=8'h03;
	15'h25ed: q<=8'h85;
	15'h25ee: q<=8'h9e;
	15'h25ef: q<=8'hbd;
	15'h25f0: q<=8'h83;
	15'h25f1: q<=8'h02;
	15'h25f2: q<=8'h30;
	15'h25f3: q<=8'h0e;
	15'h25f4: q<=8'hbc;
	15'h25f5: q<=8'hb9;
	15'h25f6: q<=8'h02;
	15'h25f7: q<=8'ha6;
	15'h25f8: q<=8'h55;
	15'h25f9: q<=8'hbd;
	15'h25fa: q<=8'h0b;
	15'h25fb: q<=8'hb6;
	15'h25fc: q<=8'h20;
	15'h25fd: q<=8'ha0;
	15'h25fe: q<=8'hbd;
	15'h25ff: q<=8'hb8;
	15'h2600: q<=8'h50;
	15'h2601: q<=8'h08;
	15'h2602: q<=8'h20;
	15'h2603: q<=8'h34;
	15'h2604: q<=8'hb6;
	15'h2605: q<=8'ha0;
	15'h2606: q<=8'h00;
	15'h2607: q<=8'h20;
	15'h2608: q<=8'hcb;
	15'h2609: q<=8'hbd;
	15'h260a: q<=8'h60;
	15'h260b: q<=8'h00;
	15'h260c: q<=8'h00;
	15'h260d: q<=8'h00;
	15'h260e: q<=8'h00;
	15'h260f: q<=8'hbd;
	15'h2610: q<=8'h8a;
	15'h2611: q<=8'h02;
	15'h2612: q<=8'h29;
	15'h2613: q<=8'h03;
	15'h2614: q<=8'ha8;
	15'h2615: q<=8'hb9;
	15'h2616: q<=8'h1e;
	15'h2617: q<=8'hb6;
	15'h2618: q<=8'hbc;
	15'h2619: q<=8'hb9;
	15'h261a: q<=8'h02;
	15'h261b: q<=8'h4c;
	15'h261c: q<=8'hfd;
	15'h261d: q<=8'hbc;
	15'h261e: q<=8'h1a;
	15'h261f: q<=8'h1a;
	15'h2620: q<=8'h4a;
	15'h2621: q<=8'h4c;
	15'h2622: q<=8'hbc;
	15'h2623: q<=8'hb9;
	15'h2624: q<=8'h02;
	15'h2625: q<=8'ha5;
	15'h2626: q<=8'h03;
	15'h2627: q<=8'h29;
	15'h2628: q<=8'h03;
	15'h2629: q<=8'h0a;
	15'h262a: q<=8'h18;
	15'h262b: q<=8'h69;
	15'h262c: q<=8'h12;
	15'h262d: q<=8'h4c;
	15'h262e: q<=8'hfd;
	15'h262f: q<=8'hbc;
	15'h2630: q<=8'h12;
	15'h2631: q<=8'h14;
	15'h2632: q<=8'h16;
	15'h2633: q<=8'h18;
	15'h2634: q<=8'ha5;
	15'h2635: q<=8'h57;
	15'h2636: q<=8'h85;
	15'h2637: q<=8'h2f;
	15'h2638: q<=8'hbc;
	15'h2639: q<=8'hb9;
	15'h263a: q<=8'h02;
	15'h263b: q<=8'hb9;
	15'h263c: q<=8'hce;
	15'h263d: q<=8'h03;
	15'h263e: q<=8'h85;
	15'h263f: q<=8'h56;
	15'h2640: q<=8'hb9;
	15'h2641: q<=8'hde;
	15'h2642: q<=8'h03;
	15'h2643: q<=8'h85;
	15'h2644: q<=8'h58;
	15'h2645: q<=8'hbd;
	15'h2646: q<=8'hcc;
	15'h2647: q<=8'h02;
	15'h2648: q<=8'h29;
	15'h2649: q<=8'h0f;
	15'h264a: q<=8'ha8;
	15'h264b: q<=8'ha5;
	15'h264c: q<=8'h56;
	15'h264d: q<=8'h49;
	15'h264e: q<=8'h80;
	15'h264f: q<=8'h18;
	15'h2650: q<=8'h79;
	15'h2651: q<=8'h8b;
	15'h2652: q<=8'hb6;
	15'h2653: q<=8'h50;
	15'h2654: q<=8'h09;
	15'h2655: q<=8'h10;
	15'h2656: q<=8'h05;
	15'h2657: q<=8'ha9;
	15'h2658: q<=8'h7f;
	15'h2659: q<=8'hb8;
	15'h265a: q<=8'h50;
	15'h265b: q<=8'h02;
	15'h265c: q<=8'ha9;
	15'h265d: q<=8'h80;
	15'h265e: q<=8'h49;
	15'h265f: q<=8'h80;
	15'h2660: q<=8'h85;
	15'h2661: q<=8'h2e;
	15'h2662: q<=8'ha5;
	15'h2663: q<=8'h58;
	15'h2664: q<=8'h49;
	15'h2665: q<=8'h80;
	15'h2666: q<=8'h18;
	15'h2667: q<=8'h79;
	15'h2668: q<=8'h87;
	15'h2669: q<=8'hb6;
	15'h266a: q<=8'h50;
	15'h266b: q<=8'h09;
	15'h266c: q<=8'h10;
	15'h266d: q<=8'h05;
	15'h266e: q<=8'ha9;
	15'h266f: q<=8'h7f;
	15'h2670: q<=8'hb8;
	15'h2671: q<=8'h50;
	15'h2672: q<=8'h02;
	15'h2673: q<=8'ha9;
	15'h2674: q<=8'h80;
	15'h2675: q<=8'h49;
	15'h2676: q<=8'h80;
	15'h2677: q<=8'h85;
	15'h2678: q<=8'h30;
	15'h2679: q<=8'hac;
	15'h267a: q<=8'h12;
	15'h267b: q<=8'h01;
	15'h267c: q<=8'hb9;
	15'h267d: q<=8'hdc;
	15'h267e: q<=8'hbc;
	15'h267f: q<=8'h85;
	15'h2680: q<=8'h59;
	15'h2681: q<=8'hb9;
	15'h2682: q<=8'hec;
	15'h2683: q<=8'hbc;
	15'h2684: q<=8'h85;
	15'h2685: q<=8'h5a;
	15'h2686: q<=8'h60;
	15'h2687: q<=8'h00;
	15'h2688: q<=8'h10;
	15'h2689: q<=8'h1f;
	15'h268a: q<=8'h28;
	15'h268b: q<=8'h2c;
	15'h268c: q<=8'h28;
	15'h268d: q<=8'h1f;
	15'h268e: q<=8'h10;
	15'h268f: q<=8'h00;
	15'h2690: q<=8'hf0;
	15'h2691: q<=8'he1;
	15'h2692: q<=8'hd8;
	15'h2693: q<=8'hd4;
	15'h2694: q<=8'hd8;
	15'h2695: q<=8'he1;
	15'h2696: q<=8'hf0;
	15'h2697: q<=8'h00;
	15'h2698: q<=8'h10;
	15'h2699: q<=8'h1f;
	15'h269a: q<=8'h28;
	15'h269b: q<=8'hbd;
	15'h269c: q<=8'hdf;
	15'h269d: q<=8'h02;
	15'h269e: q<=8'h85;
	15'h269f: q<=8'h57;
	15'h26a0: q<=8'hbc;
	15'h26a1: q<=8'hb9;
	15'h26a2: q<=8'h02;
	15'h26a3: q<=8'hb9;
	15'h26a4: q<=8'hce;
	15'h26a5: q<=8'h03;
	15'h26a6: q<=8'h85;
	15'h26a7: q<=8'h56;
	15'h26a8: q<=8'hb9;
	15'h26a9: q<=8'hde;
	15'h26aa: q<=8'h03;
	15'h26ab: q<=8'h85;
	15'h26ac: q<=8'h58;
	15'h26ad: q<=8'hbd;
	15'h26ae: q<=8'hcc;
	15'h26af: q<=8'h02;
	15'h26b0: q<=8'h10;
	15'h26b1: q<=8'h23;
	15'h26b2: q<=8'h98;
	15'h26b3: q<=8'h18;
	15'h26b4: q<=8'h69;
	15'h26b5: q<=8'h01;
	15'h26b6: q<=8'h29;
	15'h26b7: q<=8'h0f;
	15'h26b8: q<=8'ha8;
	15'h26b9: q<=8'hb9;
	15'h26ba: q<=8'hce;
	15'h26bb: q<=8'h03;
	15'h26bc: q<=8'h38;
	15'h26bd: q<=8'he5;
	15'h26be: q<=8'h56;
	15'h26bf: q<=8'h20;
	15'h26c0: q<=8'hfa;
	15'h26c1: q<=8'hb6;
	15'h26c2: q<=8'h18;
	15'h26c3: q<=8'h65;
	15'h26c4: q<=8'h56;
	15'h26c5: q<=8'h85;
	15'h26c6: q<=8'h56;
	15'h26c7: q<=8'hb9;
	15'h26c8: q<=8'hde;
	15'h26c9: q<=8'h03;
	15'h26ca: q<=8'h38;
	15'h26cb: q<=8'he5;
	15'h26cc: q<=8'h58;
	15'h26cd: q<=8'h20;
	15'h26ce: q<=8'hfa;
	15'h26cf: q<=8'hb6;
	15'h26d0: q<=8'h18;
	15'h26d1: q<=8'h65;
	15'h26d2: q<=8'h58;
	15'h26d3: q<=8'h85;
	15'h26d4: q<=8'h58;
	15'h26d5: q<=8'h20;
	15'h26d6: q<=8'h98;
	15'h26d7: q<=8'hc0;
	15'h26d8: q<=8'ha2;
	15'h26d9: q<=8'h61;
	15'h26da: q<=8'h20;
	15'h26db: q<=8'h65;
	15'h26dc: q<=8'hc7;
	15'h26dd: q<=8'ha9;
	15'h26de: q<=8'h00;
	15'h26df: q<=8'h85;
	15'h26e0: q<=8'ha9;
	15'h26e1: q<=8'h20;
	15'h26e2: q<=8'h3e;
	15'h26e3: q<=8'hbd;
	15'h26e4: q<=8'h84;
	15'h26e5: q<=8'ha9;
	15'h26e6: q<=8'ha5;
	15'h26e7: q<=8'h03;
	15'h26e8: q<=8'h29;
	15'h26e9: q<=8'h03;
	15'h26ea: q<=8'h0a;
	15'h26eb: q<=8'h18;
	15'h26ec: q<=8'h69;
	15'h26ed: q<=8'h4e;
	15'h26ee: q<=8'ha8;
	15'h26ef: q<=8'hbe;
	15'h26f0: q<=8'hc9;
	15'h26f1: q<=8'hce;
	15'h26f2: q<=8'hb9;
	15'h26f3: q<=8'hc8;
	15'h26f4: q<=8'hce;
	15'h26f5: q<=8'ha4;
	15'h26f6: q<=8'ha9;
	15'h26f7: q<=8'h4c;
	15'h26f8: q<=8'h59;
	15'h26f9: q<=8'hdf;
	15'h26fa: q<=8'h85;
	15'h26fb: q<=8'h29;
	15'h26fc: q<=8'hbd;
	15'h26fd: q<=8'hcc;
	15'h26fe: q<=8'h02;
	15'h26ff: q<=8'h29;
	15'h2700: q<=8'h07;
	15'h2701: q<=8'h85;
	15'h2702: q<=8'h2c;
	15'h2703: q<=8'h86;
	15'h2704: q<=8'h2b;
	15'h2705: q<=8'ha2;
	15'h2706: q<=8'h02;
	15'h2707: q<=8'ha9;
	15'h2708: q<=8'h00;
	15'h2709: q<=8'h46;
	15'h270a: q<=8'h2c;
	15'h270b: q<=8'h90;
	15'h270c: q<=8'h03;
	15'h270d: q<=8'h18;
	15'h270e: q<=8'h65;
	15'h270f: q<=8'h29;
	15'h2710: q<=8'h0a;
	15'h2711: q<=8'h08;
	15'h2712: q<=8'h6a;
	15'h2713: q<=8'h28;
	15'h2714: q<=8'h6a;
	15'h2715: q<=8'hca;
	15'h2716: q<=8'h10;
	15'h2717: q<=8'hf1;
	15'h2718: q<=8'ha6;
	15'h2719: q<=8'h2b;
	15'h271a: q<=8'h60;
	15'h271b: q<=8'ha9;
	15'h271c: q<=8'h04;
	15'h271d: q<=8'hac;
	15'h271e: q<=8'h48;
	15'h271f: q<=8'h01;
	15'h2720: q<=8'h30;
	15'h2721: q<=8'h02;
	15'h2722: q<=8'ha9;
	15'h2723: q<=8'h00;
	15'h2724: q<=8'h85;
	15'h2725: q<=8'h9e;
	15'h2726: q<=8'had;
	15'h2727: q<=8'h48;
	15'h2728: q<=8'h01;
	15'h2729: q<=8'h18;
	15'h272a: q<=8'h69;
	15'h272b: q<=8'h40;
	15'h272c: q<=8'h4a;
	15'h272d: q<=8'h4a;
	15'h272e: q<=8'h4a;
	15'h272f: q<=8'h4a;
	15'h2730: q<=8'hc9;
	15'h2731: q<=8'h05;
	15'h2732: q<=8'h90;
	15'h2733: q<=8'h02;
	15'h2734: q<=8'ha9;
	15'h2735: q<=8'h00;
	15'h2736: q<=8'ha8;
	15'h2737: q<=8'hb9;
	15'h2738: q<=8'h55;
	15'h2739: q<=8'hb7;
	15'h273a: q<=8'h85;
	15'h273b: q<=8'h29;
	15'h273c: q<=8'hbd;
	15'h273d: q<=8'h83;
	15'h273e: q<=8'h02;
	15'h273f: q<=8'h30;
	15'h2740: q<=8'h0b;
	15'h2741: q<=8'hbc;
	15'h2742: q<=8'hb9;
	15'h2743: q<=8'h02;
	15'h2744: q<=8'ha5;
	15'h2745: q<=8'h29;
	15'h2746: q<=8'h20;
	15'h2747: q<=8'ha0;
	15'h2748: q<=8'hbd;
	15'h2749: q<=8'hb8;
	15'h274a: q<=8'h50;
	15'h274b: q<=8'h08;
	15'h274c: q<=8'h20;
	15'h274d: q<=8'h34;
	15'h274e: q<=8'hb6;
	15'h274f: q<=8'ha4;
	15'h2750: q<=8'h29;
	15'h2751: q<=8'h20;
	15'h2752: q<=8'hcb;
	15'h2753: q<=8'hbd;
	15'h2754: q<=8'h60;
	15'h2755: q<=8'h0d;
	15'h2756: q<=8'h0c;
	15'h2757: q<=8'h0b;
	15'h2758: q<=8'h0a;
	15'h2759: q<=8'h09;
	15'h275a: q<=8'h09;
	15'h275b: q<=8'ha2;
	15'h275c: q<=8'h0b;
	15'h275d: q<=8'h86;
	15'h275e: q<=8'h37;
	15'h275f: q<=8'ha6;
	15'h2760: q<=8'h37;
	15'h2761: q<=8'hbd;
	15'h2762: q<=8'hd3;
	15'h2763: q<=8'h02;
	15'h2764: q<=8'hf0;
	15'h2765: q<=8'h1b;
	15'h2766: q<=8'h85;
	15'h2767: q<=8'h57;
	15'h2768: q<=8'h85;
	15'h2769: q<=8'h2f;
	15'h276a: q<=8'he0;
	15'h276b: q<=8'h08;
	15'h276c: q<=8'hbc;
	15'h276d: q<=8'had;
	15'h276e: q<=8'h02;
	15'h276f: q<=8'hb0;
	15'h2770: q<=8'h05;
	15'h2771: q<=8'ha9;
	15'h2772: q<=8'h08;
	15'h2773: q<=8'hb8;
	15'h2774: q<=8'h50;
	15'h2775: q<=8'h08;
	15'h2776: q<=8'ha5;
	15'h2777: q<=8'h03;
	15'h2778: q<=8'h0a;
	15'h2779: q<=8'h29;
	15'h277a: q<=8'h06;
	15'h277b: q<=8'h18;
	15'h277c: q<=8'h69;
	15'h277d: q<=8'h20;
	15'h277e: q<=8'h20;
	15'h277f: q<=8'hfd;
	15'h2780: q<=8'hbc;
	15'h2781: q<=8'hc6;
	15'h2782: q<=8'h37;
	15'h2783: q<=8'h10;
	15'h2784: q<=8'hda;
	15'h2785: q<=8'ha0;
	15'h2786: q<=8'h04;
	15'h2787: q<=8'had;
	15'h2788: q<=8'h35;
	15'h2789: q<=8'h01;
	15'h278a: q<=8'hc9;
	15'h278b: q<=8'h06;
	15'h278c: q<=8'h90;
	15'h278d: q<=8'h08;
	15'h278e: q<=8'ha0;
	15'h278f: q<=8'h0b;
	15'h2790: q<=8'hc9;
	15'h2791: q<=8'h08;
	15'h2792: q<=8'h90;
	15'h2793: q<=8'h02;
	15'h2794: q<=8'ha0;
	15'h2795: q<=8'h0c;
	15'h2796: q<=8'h8c;
	15'h2797: q<=8'h08;
	15'h2798: q<=8'h08;
	15'h2799: q<=8'h60;
	15'h279a: q<=8'ha0;
	15'h279b: q<=8'h00;
	15'h279c: q<=8'h84;
	15'h279d: q<=8'h9e;
	15'h279e: q<=8'ha2;
	15'h279f: q<=8'h07;
	15'h27a0: q<=8'h86;
	15'h27a1: q<=8'h37;
	15'h27a2: q<=8'ha6;
	15'h27a3: q<=8'h37;
	15'h27a4: q<=8'hbd;
	15'h27a5: q<=8'h0a;
	15'h27a6: q<=8'h03;
	15'h27a7: q<=8'hf0;
	15'h27a8: q<=8'h29;
	15'h27a9: q<=8'h85;
	15'h27aa: q<=8'h57;
	15'h27ab: q<=8'hbd;
	15'h27ac: q<=8'hfa;
	15'h27ad: q<=8'h02;
	15'h27ae: q<=8'h85;
	15'h27af: q<=8'h29;
	15'h27b0: q<=8'hbc;
	15'h27b1: q<=8'h02;
	15'h27b2: q<=8'h03;
	15'h27b3: q<=8'hc0;
	15'h27b4: q<=8'h01;
	15'h27b5: q<=8'hd0;
	15'h27b6: q<=8'h06;
	15'h27b7: q<=8'h20;
	15'h27b8: q<=8'heb;
	15'h27b9: q<=8'hb7;
	15'h27ba: q<=8'hb8;
	15'h27bb: q<=8'h50;
	15'h27bc: q<=8'h15;
	15'h27bd: q<=8'hbd;
	15'h27be: q<=8'h12;
	15'h27bf: q<=8'h03;
	15'h27c0: q<=8'h4a;
	15'h27c1: q<=8'h29;
	15'h27c2: q<=8'hfe;
	15'h27c3: q<=8'hc0;
	15'h27c4: q<=8'h02;
	15'h27c5: q<=8'h90;
	15'h27c6: q<=8'h02;
	15'h27c7: q<=8'ha9;
	15'h27c8: q<=8'h00;
	15'h27c9: q<=8'h18;
	15'h27ca: q<=8'h79;
	15'h27cb: q<=8'he5;
	15'h27cc: q<=8'hb7;
	15'h27cd: q<=8'ha4;
	15'h27ce: q<=8'h29;
	15'h27cf: q<=8'h20;
	15'h27d0: q<=8'hfd;
	15'h27d1: q<=8'hbc;
	15'h27d2: q<=8'hc6;
	15'h27d3: q<=8'h37;
	15'h27d4: q<=8'h10;
	15'h27d5: q<=8'hcc;
	15'h27d6: q<=8'had;
	15'h27d7: q<=8'h20;
	15'h27d8: q<=8'h07;
	15'h27d9: q<=8'hf0;
	15'h27da: q<=8'h09;
	15'h27db: q<=8'ha5;
	15'h27dc: q<=8'h9f;
	15'h27dd: q<=8'hc9;
	15'h27de: q<=8'h0d;
	15'h27df: q<=8'h90;
	15'h27e0: q<=8'h03;
	15'h27e1: q<=8'h8d;
	15'h27e2: q<=8'hff;
	15'h27e3: q<=8'h01;
	15'h27e4: q<=8'h60;
	15'h27e5: q<=8'h00;
	15'h27e6: q<=8'h00;
	15'h27e7: q<=8'h5a;
	15'h27e8: q<=8'h58;
	15'h27e9: q<=8'h56;
	15'h27ea: q<=8'h1c;
	15'h27eb: q<=8'ha4;
	15'h27ec: q<=8'h29;
	15'h27ed: q<=8'hb9;
	15'h27ee: q<=8'h35;
	15'h27ef: q<=8'h04;
	15'h27f0: q<=8'h85;
	15'h27f1: q<=8'h56;
	15'h27f2: q<=8'hb9;
	15'h27f3: q<=8'h45;
	15'h27f4: q<=8'h04;
	15'h27f5: q<=8'h85;
	15'h27f6: q<=8'h58;
	15'h27f7: q<=8'h20;
	15'h27f8: q<=8'h98;
	15'h27f9: q<=8'hc0;
	15'h27fa: q<=8'ha2;
	15'h27fb: q<=8'h61;
	15'h27fc: q<=8'h20;
	15'h27fd: q<=8'h65;
	15'h27fe: q<=8'hc7;
	15'h27ff: q<=8'hae;
	15'h2800: q<=8'h3b;
	15'h2801: q<=8'h01;
	15'h2802: q<=8'hce;
	15'h2803: q<=8'h3c;
	15'h2804: q<=8'h01;
	15'h2805: q<=8'hd0;
	15'h2806: q<=8'h0a;
	15'h2807: q<=8'he8;
	15'h2808: q<=8'h8e;
	15'h2809: q<=8'h3b;
	15'h280a: q<=8'h01;
	15'h280b: q<=8'hbd;
	15'h280c: q<=8'h2a;
	15'h280d: q<=8'hb8;
	15'h280e: q<=8'h8d;
	15'h280f: q<=8'h3c;
	15'h2810: q<=8'h01;
	15'h2811: q<=8'hbc;
	15'h2812: q<=8'h3d;
	15'h2813: q<=8'hb8;
	15'h2814: q<=8'h30;
	15'h2815: q<=8'h03;
	15'h2816: q<=8'h20;
	15'h2817: q<=8'h4e;
	15'h2818: q<=8'hb8;
	15'h2819: q<=8'had;
	15'h281a: q<=8'h3b;
	15'h281b: q<=8'h01;
	15'h281c: q<=8'h0a;
	15'h281d: q<=8'h18;
	15'h281e: q<=8'h69;
	15'h281f: q<=8'h28;
	15'h2820: q<=8'ha8;
	15'h2821: q<=8'hbe;
	15'h2822: q<=8'hc9;
	15'h2823: q<=8'hce;
	15'h2824: q<=8'hb9;
	15'h2825: q<=8'hc8;
	15'h2826: q<=8'hce;
	15'h2827: q<=8'h4c;
	15'h2828: q<=8'h57;
	15'h2829: q<=8'hdf;
	15'h282a: q<=8'h02;
	15'h282b: q<=8'h02;
	15'h282c: q<=8'h02;
	15'h282d: q<=8'h02;
	15'h282e: q<=8'h02;
	15'h282f: q<=8'h04;
	15'h2830: q<=8'h03;
	15'h2831: q<=8'h02;
	15'h2832: q<=8'h01;
	15'h2833: q<=8'h20;
	15'h2834: q<=8'h03;
	15'h2835: q<=8'h03;
	15'h2836: q<=8'h03;
	15'h2837: q<=8'h03;
	15'h2838: q<=8'h03;
	15'h2839: q<=8'h03;
	15'h283a: q<=8'h03;
	15'h283b: q<=8'h3b;
	15'h283c: q<=8'hb8;
	15'h283d: q<=8'h00;
	15'h283e: q<=8'h02;
	15'h283f: q<=8'h02;
	15'h2840: q<=8'h02;
	15'h2841: q<=8'h02;
	15'h2842: q<=8'h02;
	15'h2843: q<=8'h02;
	15'h2844: q<=8'h02;
	15'h2845: q<=8'h04;
	15'h2846: q<=8'h06;
	15'h2847: q<=8'hff;
	15'h2848: q<=8'hff;
	15'h2849: q<=8'hff;
	15'h284a: q<=8'hff;
	15'h284b: q<=8'hff;
	15'h284c: q<=8'hff;
	15'h284d: q<=8'hff;
	15'h284e: q<=8'hb9;
	15'h284f: q<=8'h58;
	15'h2850: q<=8'hb8;
	15'h2851: q<=8'h48;
	15'h2852: q<=8'hb9;
	15'h2853: q<=8'h57;
	15'h2854: q<=8'hb8;
	15'h2855: q<=8'h48;
	15'h2856: q<=8'h60;
	15'h2857: q<=8'h5e;
	15'h2858: q<=8'hb8;
	15'h2859: q<=8'h74;
	15'h285a: q<=8'hb8;
	15'h285b: q<=8'h87;
	15'h285c: q<=8'hb8;
	15'h285d: q<=8'h95;
	15'h285e: q<=8'hb8;
	15'h285f: q<=8'ha9;
	15'h2860: q<=8'h0c;
	15'h2861: q<=8'h8d;
	15'h2862: q<=8'h0b;
	15'h2863: q<=8'h08;
	15'h2864: q<=8'h85;
	15'h2865: q<=8'h24;
	15'h2866: q<=8'ha9;
	15'h2867: q<=8'h04;
	15'h2868: q<=8'h8d;
	15'h2869: q<=8'h0a;
	15'h286a: q<=8'h08;
	15'h286b: q<=8'h85;
	15'h286c: q<=8'h23;
	15'h286d: q<=8'ha9;
	15'h286e: q<=8'h00;
	15'h286f: q<=8'h85;
	15'h2870: q<=8'h22;
	15'h2871: q<=8'h8d;
	15'h2872: q<=8'h09;
	15'h2873: q<=8'h08;
	15'h2874: q<=8'h60;
	15'h2875: q<=8'ha4;
	15'h2876: q<=8'h22;
	15'h2877: q<=8'ha2;
	15'h2878: q<=8'h02;
	15'h2879: q<=8'hb5;
	15'h287a: q<=8'h22;
	15'h287b: q<=8'h48;
	15'h287c: q<=8'h94;
	15'h287d: q<=8'h22;
	15'h287e: q<=8'h98;
	15'h287f: q<=8'h9d;
	15'h2880: q<=8'h09;
	15'h2881: q<=8'h08;
	15'h2882: q<=8'h68;
	15'h2883: q<=8'ha8;
	15'h2884: q<=8'hca;
	15'h2885: q<=8'h10;
	15'h2886: q<=8'hf2;
	15'h2887: q<=8'h60;
	15'h2888: q<=8'h20;
	15'h2889: q<=8'h96;
	15'h288a: q<=8'hc1;
	15'h288b: q<=8'ha9;
	15'h288c: q<=8'h7f;
	15'h288d: q<=8'h8d;
	15'h288e: q<=8'h39;
	15'h288f: q<=8'h01;
	15'h2890: q<=8'ha9;
	15'h2891: q<=8'h04;
	15'h2892: q<=8'h8d;
	15'h2893: q<=8'h3a;
	15'h2894: q<=8'h01;
	15'h2895: q<=8'h60;
	15'h2896: q<=8'had;
	15'h2897: q<=8'h39;
	15'h2898: q<=8'h01;
	15'h2899: q<=8'h8d;
	15'h289a: q<=8'hfc;
	15'h289b: q<=8'h2f;
	15'h289c: q<=8'had;
	15'h289d: q<=8'h3a;
	15'h289e: q<=8'h01;
	15'h289f: q<=8'h09;
	15'h28a0: q<=8'h70;
	15'h28a1: q<=8'h8d;
	15'h28a2: q<=8'hfd;
	15'h28a3: q<=8'h2f;
	15'h28a4: q<=8'ha9;
	15'h28a5: q<=8'hc0;
	15'h28a6: q<=8'h8d;
	15'h28a7: q<=8'hff;
	15'h28a8: q<=8'h2f;
	15'h28a9: q<=8'had;
	15'h28aa: q<=8'h39;
	15'h28ab: q<=8'h01;
	15'h28ac: q<=8'h38;
	15'h28ad: q<=8'he9;
	15'h28ae: q<=8'h20;
	15'h28af: q<=8'h10;
	15'h28b0: q<=8'h05;
	15'h28b1: q<=8'h29;
	15'h28b2: q<=8'h7f;
	15'h28b3: q<=8'hce;
	15'h28b4: q<=8'h3a;
	15'h28b5: q<=8'h01;
	15'h28b6: q<=8'h8d;
	15'h28b7: q<=8'h39;
	15'h28b8: q<=8'h01;
	15'h28b9: q<=8'h60;
	15'h28ba: q<=8'ha9;
	15'h28bb: q<=8'h3f;
	15'h28bc: q<=8'ha2;
	15'h28bd: q<=8'hf2;
	15'h28be: q<=8'h20;
	15'h28bf: q<=8'h39;
	15'h28c0: q<=8'hdf;
	15'h28c1: q<=8'ha9;
	15'h28c2: q<=8'h00;
	15'h28c3: q<=8'h85;
	15'h28c4: q<=8'h6a;
	15'h28c5: q<=8'h85;
	15'h28c6: q<=8'h6b;
	15'h28c7: q<=8'h85;
	15'h28c8: q<=8'h6c;
	15'h28c9: q<=8'h85;
	15'h28ca: q<=8'h6d;
	15'h28cb: q<=8'h8d;
	15'h28cc: q<=8'h02;
	15'h28cd: q<=8'h02;
	15'h28ce: q<=8'h85;
	15'h28cf: q<=8'h68;
	15'h28d0: q<=8'h85;
	15'h28d1: q<=8'h69;
	15'h28d2: q<=8'ha9;
	15'h28d3: q<=8'he0;
	15'h28d4: q<=8'h85;
	15'h28d5: q<=8'h5f;
	15'h28d6: q<=8'ha9;
	15'h28d7: q<=8'hff;
	15'h28d8: q<=8'h85;
	15'h28d9: q<=8'h5b;
	15'h28da: q<=8'h20;
	15'h28db: q<=8'h67;
	15'h28dc: q<=8'hb9;
	15'h28dd: q<=8'h85;
	15'h28de: q<=8'h77;
	15'h28df: q<=8'h86;
	15'h28e0: q<=8'h76;
	15'h28e1: q<=8'ha2;
	15'h28e2: q<=8'h0f;
	15'h28e3: q<=8'h86;
	15'h28e4: q<=8'h37;
	15'h28e5: q<=8'ha6;
	15'h28e6: q<=8'h37;
	15'h28e7: q<=8'hbd;
	15'h28e8: q<=8'h83;
	15'h28e9: q<=8'h02;
	15'h28ea: q<=8'hf0;
	15'h28eb: q<=8'h49;
	15'h28ec: q<=8'h85;
	15'h28ed: q<=8'h57;
	15'h28ee: q<=8'hbd;
	15'h28ef: q<=8'h63;
	15'h28f0: q<=8'h02;
	15'h28f1: q<=8'h85;
	15'h28f2: q<=8'h56;
	15'h28f3: q<=8'hbd;
	15'h28f4: q<=8'ha3;
	15'h28f5: q<=8'h02;
	15'h28f6: q<=8'h85;
	15'h28f7: q<=8'h58;
	15'h28f8: q<=8'h20;
	15'h28f9: q<=8'h98;
	15'h28fa: q<=8'hc0;
	15'h28fb: q<=8'ha9;
	15'h28fc: q<=8'h00;
	15'h28fd: q<=8'h85;
	15'h28fe: q<=8'h73;
	15'h28ff: q<=8'h20;
	15'h2900: q<=8'h44;
	15'h2901: q<=8'hb9;
	15'h2902: q<=8'h20;
	15'h2903: q<=8'hba;
	15'h2904: q<=8'hc3;
	15'h2905: q<=8'ha9;
	15'h2906: q<=8'ha0;
	15'h2907: q<=8'h20;
	15'h2908: q<=8'h6a;
	15'h2909: q<=8'hb5;
	15'h290a: q<=8'h20;
	15'h290b: q<=8'h44;
	15'h290c: q<=8'hb9;
	15'h290d: q<=8'ha2;
	15'h290e: q<=8'h61;
	15'h290f: q<=8'h20;
	15'h2910: q<=8'h72;
	15'h2911: q<=8'hc7;
	15'h2912: q<=8'h20;
	15'h2913: q<=8'h55;
	15'h2914: q<=8'hb9;
	15'h2915: q<=8'h20;
	15'h2916: q<=8'h6c;
	15'h2917: q<=8'hdf;
	15'h2918: q<=8'ha5;
	15'h2919: q<=8'h37;
	15'h291a: q<=8'h29;
	15'h291b: q<=8'h07;
	15'h291c: q<=8'hc9;
	15'h291d: q<=8'h07;
	15'h291e: q<=8'hd0;
	15'h291f: q<=8'h02;
	15'h2920: q<=8'ha9;
	15'h2921: q<=8'h00;
	15'h2922: q<=8'ha8;
	15'h2923: q<=8'h84;
	15'h2924: q<=8'h9e;
	15'h2925: q<=8'ha9;
	15'h2926: q<=8'h08;
	15'h2927: q<=8'h20;
	15'h2928: q<=8'h4c;
	15'h2929: q<=8'hdf;
	15'h292a: q<=8'ha9;
	15'h292b: q<=8'h00;
	15'h292c: q<=8'h20;
	15'h292d: q<=8'h4a;
	15'h292e: q<=8'hdf;
	15'h292f: q<=8'h20;
	15'h2930: q<=8'h67;
	15'h2931: q<=8'hb9;
	15'h2932: q<=8'h20;
	15'h2933: q<=8'h39;
	15'h2934: q<=8'hdf;
	15'h2935: q<=8'hc6;
	15'h2936: q<=8'h37;
	15'h2937: q<=8'h10;
	15'h2938: q<=8'hac;
	15'h2939: q<=8'h20;
	15'h293a: q<=8'h44;
	15'h293b: q<=8'hb9;
	15'h293c: q<=8'ha9;
	15'h293d: q<=8'h01;
	15'h293e: q<=8'h20;
	15'h293f: q<=8'h6a;
	15'h2940: q<=8'hdf;
	15'h2941: q<=8'h20;
	15'h2942: q<=8'h09;
	15'h2943: q<=8'hdf;
	15'h2944: q<=8'ha6;
	15'h2945: q<=8'h74;
	15'h2946: q<=8'ha4;
	15'h2947: q<=8'h75;
	15'h2948: q<=8'ha5;
	15'h2949: q<=8'h76;
	15'h294a: q<=8'h85;
	15'h294b: q<=8'h74;
	15'h294c: q<=8'h86;
	15'h294d: q<=8'h76;
	15'h294e: q<=8'ha5;
	15'h294f: q<=8'h77;
	15'h2950: q<=8'h85;
	15'h2951: q<=8'h75;
	15'h2952: q<=8'h84;
	15'h2953: q<=8'h77;
	15'h2954: q<=8'h60;
	15'h2955: q<=8'ha5;
	15'h2956: q<=8'h57;
	15'h2957: q<=8'h4a;
	15'h2958: q<=8'h4a;
	15'h2959: q<=8'h4a;
	15'h295a: q<=8'h4a;
	15'h295b: q<=8'ha0;
	15'h295c: q<=8'h00;
	15'h295d: q<=8'hc8;
	15'h295e: q<=8'h4a;
	15'h295f: q<=8'hd0;
	15'h2960: q<=8'hfc;
	15'h2961: q<=8'h18;
	15'h2962: q<=8'h69;
	15'h2963: q<=8'h02;
	15'h2964: q<=8'ha0;
	15'h2965: q<=8'h00;
	15'h2966: q<=8'h60;
	15'h2967: q<=8'had;
	15'h2968: q<=8'h15;
	15'h2969: q<=8'h04;
	15'h296a: q<=8'hf0;
	15'h296b: q<=8'h09;
	15'h296c: q<=8'had;
	15'h296d: q<=8'h6f;
	15'h296e: q<=8'hce;
	15'h296f: q<=8'hae;
	15'h2970: q<=8'h6e;
	15'h2971: q<=8'hce;
	15'h2972: q<=8'hb8;
	15'h2973: q<=8'h50;
	15'h2974: q<=8'h06;
	15'h2975: q<=8'had;
	15'h2976: q<=8'h87;
	15'h2977: q<=8'hce;
	15'h2978: q<=8'hae;
	15'h2979: q<=8'h86;
	15'h297a: q<=8'hce;
	15'h297b: q<=8'h60;
	15'h297c: q<=8'hf0;
	15'h297d: q<=8'he7;
	15'h297e: q<=8'hcf;
	15'h297f: q<=8'haa;
	15'h2980: q<=8'h80;
	15'h2981: q<=8'h56;
	15'h2982: q<=8'h31;
	15'h2983: q<=8'h19;
	15'h2984: q<=8'h10;
	15'h2985: q<=8'h19;
	15'h2986: q<=8'h31;
	15'h2987: q<=8'h56;
	15'h2988: q<=8'h80;
	15'h2989: q<=8'haa;
	15'h298a: q<=8'hcf;
	15'h298b: q<=8'he7;
	15'h298c: q<=8'hf0;
	15'h298d: q<=8'hf0;
	15'h298e: q<=8'hf0;
	15'h298f: q<=8'hb8;
	15'h2990: q<=8'h80;
	15'h2991: q<=8'h48;
	15'h2992: q<=8'h10;
	15'h2993: q<=8'h10;
	15'h2994: q<=8'h10;
	15'h2995: q<=8'h10;
	15'h2996: q<=8'h10;
	15'h2997: q<=8'h48;
	15'h2998: q<=8'h80;
	15'h2999: q<=8'hb8;
	15'h299a: q<=8'hf0;
	15'h299b: q<=8'hf0;
	15'h299c: q<=8'hf0;
	15'h299d: q<=8'hf0;
	15'h299e: q<=8'hb8;
	15'h299f: q<=8'hb8;
	15'h29a0: q<=8'h80;
	15'h29a1: q<=8'h48;
	15'h29a2: q<=8'h48;
	15'h29a3: q<=8'h10;
	15'h29a4: q<=8'h10;
	15'h29a5: q<=8'h10;
	15'h29a6: q<=8'h48;
	15'h29a7: q<=8'h48;
	15'h29a8: q<=8'h80;
	15'h29a9: q<=8'hb8;
	15'h29aa: q<=8'hb8;
	15'h29ab: q<=8'hf0;
	15'h29ac: q<=8'hec;
	15'h29ad: q<=8'hd5;
	15'h29ae: q<=8'hb1;
	15'h29af: q<=8'h90;
	15'h29b0: q<=8'h70;
	15'h29b1: q<=8'h4f;
	15'h29b2: q<=8'h2b;
	15'h29b3: q<=8'h14;
	15'h29b4: q<=8'h14;
	15'h29b5: q<=8'h2b;
	15'h29b6: q<=8'h4f;
	15'h29b7: q<=8'h70;
	15'h29b8: q<=8'h90;
	15'h29b9: q<=8'hb1;
	15'h29ba: q<=8'hd5;
	15'h29bb: q<=8'hec;
	15'h29bc: q<=8'hf0;
	15'h29bd: q<=8'hc0;
	15'h29be: q<=8'ha0;
	15'h29bf: q<=8'h94;
	15'h29c0: q<=8'h6c;
	15'h29c1: q<=8'h60;
	15'h29c2: q<=8'h40;
	15'h29c3: q<=8'h10;
	15'h29c4: q<=8'h10;
	15'h29c5: q<=8'h40;
	15'h29c6: q<=8'h60;
	15'h29c7: q<=8'h6c;
	15'h29c8: q<=8'h94;
	15'h29c9: q<=8'ha0;
	15'h29ca: q<=8'hc0;
	15'h29cb: q<=8'hf0;
	15'h29cc: q<=8'hd9;
	15'h29cd: q<=8'hc2;
	15'h29ce: q<=8'hac;
	15'h29cf: q<=8'h97;
	15'h29d0: q<=8'h80;
	15'h29d1: q<=8'h69;
	15'h29d2: q<=8'h52;
	15'h29d3: q<=8'h3c;
	15'h29d4: q<=8'h27;
	15'h29d5: q<=8'h10;
	15'h29d6: q<=8'h35;
	15'h29d7: q<=8'h5a;
	15'h29d8: q<=8'h80;
	15'h29d9: q<=8'ha6;
	15'h29da: q<=8'hca;
	15'h29db: q<=8'hf0;
	15'h29dc: q<=8'hea;
	15'h29dd: q<=8'he0;
	15'h29de: q<=8'h9c;
	15'h29df: q<=8'h80;
	15'h29e0: q<=8'h64;
	15'h29e1: q<=8'h20;
	15'h29e2: q<=8'h16;
	15'h29e3: q<=8'h50;
	15'h29e4: q<=8'h16;
	15'h29e5: q<=8'h20;
	15'h29e6: q<=8'h64;
	15'h29e7: q<=8'h80;
	15'h29e8: q<=8'h9c;
	15'h29e9: q<=8'he0;
	15'h29ea: q<=8'hea;
	15'h29eb: q<=8'hb0;
	15'h29ec: q<=8'h10;
	15'h29ed: q<=8'h1e;
	15'h29ee: q<=8'h2c;
	15'h29ef: q<=8'h3a;
	15'h29f0: q<=8'h48;
	15'h29f1: q<=8'h56;
	15'h29f2: q<=8'h64;
	15'h29f3: q<=8'h70;
	15'h29f4: q<=8'h90;
	15'h29f5: q<=8'h9e;
	15'h29f6: q<=8'hac;
	15'h29f7: q<=8'hba;
	15'h29f8: q<=8'hc8;
	15'h29f9: q<=8'hd6;
	15'h29fa: q<=8'he4;
	15'h29fb: q<=8'hf0;
	15'h29fc: q<=8'h10;
	15'h29fd: q<=8'h1e;
	15'h29fe: q<=8'h2d;
	15'h29ff: q<=8'h3c;
	15'h2a00: q<=8'h4b;
	15'h2a01: q<=8'h5a;
	15'h2a02: q<=8'h69;
	15'h2a03: q<=8'h78;
	15'h2a04: q<=8'h87;
	15'h2a05: q<=8'h96;
	15'h2a06: q<=8'ha5;
	15'h2a07: q<=8'hb4;
	15'h2a08: q<=8'hc3;
	15'h2a09: q<=8'hd2;
	15'h2a0a: q<=8'he1;
	15'h2a0b: q<=8'hf0;
	15'h2a0c: q<=8'h10;
	15'h2a0d: q<=8'h10;
	15'h2a0e: q<=8'h10;
	15'h2a0f: q<=8'h10;
	15'h2a10: q<=8'h16;
	15'h2a11: q<=8'h29;
	15'h2a12: q<=8'h46;
	15'h2a13: q<=8'h69;
	15'h2a14: q<=8'h97;
	15'h2a15: q<=8'hba;
	15'h2a16: q<=8'hd7;
	15'h2a17: q<=8'hea;
	15'h2a18: q<=8'hf0;
	15'h2a19: q<=8'hf0;
	15'h2a1a: q<=8'hf0;
	15'h2a1b: q<=8'hf0;
	15'h2a1c: q<=8'h10;
	15'h2a1d: q<=8'h24;
	15'h2a1e: q<=8'h30;
	15'h2a1f: q<=8'h36;
	15'h2a20: q<=8'h3e;
	15'h2a21: q<=8'h49;
	15'h2a22: q<=8'h5a;
	15'h2a23: q<=8'h75;
	15'h2a24: q<=8'h94;
	15'h2a25: q<=8'ha4;
	15'h2a26: q<=8'hac;
	15'h2a27: q<=8'hba;
	15'h2a28: q<=8'hda;
	15'h2a29: q<=8'he2;
	15'h2a2a: q<=8'hea;
	15'h2a2b: q<=8'hf0;
	15'h2a2c: q<=8'h80;
	15'h2a2d: q<=8'h70;
	15'h2a2e: q<=8'h48;
	15'h2a2f: q<=8'h20;
	15'h2a30: q<=8'h10;
	15'h2a31: q<=8'h20;
	15'h2a32: q<=8'h48;
	15'h2a33: q<=8'h70;
	15'h2a34: q<=8'h80;
	15'h2a35: q<=8'h90;
	15'h2a36: q<=8'hb8;
	15'h2a37: q<=8'he0;
	15'h2a38: q<=8'hf0;
	15'h2a39: q<=8'he0;
	15'h2a3a: q<=8'hb8;
	15'h2a3b: q<=8'h90;
	15'h2a3c: q<=8'hda;
	15'h2a3d: q<=8'ha4;
	15'h2a3e: q<=8'h87;
	15'h2a3f: q<=8'h80;
	15'h2a40: q<=8'h79;
	15'h2a41: q<=8'h5c;
	15'h2a42: q<=8'h26;
	15'h2a43: q<=8'h10;
	15'h2a44: q<=8'h10;
	15'h2a45: q<=8'h20;
	15'h2a46: q<=8'h48;
	15'h2a47: q<=8'h80;
	15'h2a48: q<=8'hb8;
	15'h2a49: q<=8'he0;
	15'h2a4a: q<=8'hf0;
	15'h2a4b: q<=8'hf0;
	15'h2a4c: q<=8'h10;
	15'h2a4d: q<=8'h10;
	15'h2a4e: q<=8'h30;
	15'h2a4f: q<=8'h30;
	15'h2a50: q<=8'h50;
	15'h2a51: q<=8'h50;
	15'h2a52: q<=8'h70;
	15'h2a53: q<=8'h70;
	15'h2a54: q<=8'h90;
	15'h2a55: q<=8'h90;
	15'h2a56: q<=8'hb0;
	15'h2a57: q<=8'hb0;
	15'h2a58: q<=8'hd0;
	15'h2a59: q<=8'hd0;
	15'h2a5a: q<=8'hf0;
	15'h2a5b: q<=8'hf0;
	15'h2a5c: q<=8'hb0;
	15'h2a5d: q<=8'h80;
	15'h2a5e: q<=8'h50;
	15'h2a5f: q<=8'h47;
	15'h2a60: q<=8'h18;
	15'h2a61: q<=8'h30;
	15'h2a62: q<=8'h18;
	15'h2a63: q<=8'h47;
	15'h2a64: q<=8'h50;
	15'h2a65: q<=8'h80;
	15'h2a66: q<=8'hb0;
	15'h2a67: q<=8'hb9;
	15'h2a68: q<=8'he8;
	15'h2a69: q<=8'hd4;
	15'h2a6a: q<=8'he8;
	15'h2a6b: q<=8'hb9;
	15'h2a6c: q<=8'h10;
	15'h2a6d: q<=8'h1e;
	15'h2a6e: q<=8'h21;
	15'h2a6f: q<=8'h28;
	15'h2a70: q<=8'h3c;
	15'h2a71: q<=8'h55;
	15'h2a72: q<=8'h66;
	15'h2a73: q<=8'h73;
	15'h2a74: q<=8'h8d;
	15'h2a75: q<=8'h9a;
	15'h2a76: q<=8'hab;
	15'h2a77: q<=8'hc4;
	15'h2a78: q<=8'hd8;
	15'h2a79: q<=8'hdf;
	15'h2a7a: q<=8'he2;
	15'h2a7b: q<=8'hf0;
	15'h2a7c: q<=8'h80;
	15'h2a7d: q<=8'haa;
	15'h2a7e: q<=8'hcf;
	15'h2a7f: q<=8'he7;
	15'h2a80: q<=8'hf0;
	15'h2a81: q<=8'he7;
	15'h2a82: q<=8'hcf;
	15'h2a83: q<=8'haa;
	15'h2a84: q<=8'h80;
	15'h2a85: q<=8'h56;
	15'h2a86: q<=8'h31;
	15'h2a87: q<=8'h19;
	15'h2a88: q<=8'h10;
	15'h2a89: q<=8'h19;
	15'h2a8a: q<=8'h31;
	15'h2a8b: q<=8'h56;
	15'h2a8c: q<=8'h80;
	15'h2a8d: q<=8'hb8;
	15'h2a8e: q<=8'hf0;
	15'h2a8f: q<=8'hf0;
	15'h2a90: q<=8'hf0;
	15'h2a91: q<=8'hf0;
	15'h2a92: q<=8'hf0;
	15'h2a93: q<=8'hb8;
	15'h2a94: q<=8'h80;
	15'h2a95: q<=8'h48;
	15'h2a96: q<=8'h10;
	15'h2a97: q<=8'h10;
	15'h2a98: q<=8'h10;
	15'h2a99: q<=8'h10;
	15'h2a9a: q<=8'h10;
	15'h2a9b: q<=8'h48;
	15'h2a9c: q<=8'h80;
	15'h2a9d: q<=8'hb8;
	15'h2a9e: q<=8'hb8;
	15'h2a9f: q<=8'hf0;
	15'h2aa0: q<=8'hf0;
	15'h2aa1: q<=8'hf0;
	15'h2aa2: q<=8'hb8;
	15'h2aa3: q<=8'hb8;
	15'h2aa4: q<=8'h80;
	15'h2aa5: q<=8'h48;
	15'h2aa6: q<=8'h48;
	15'h2aa7: q<=8'h10;
	15'h2aa8: q<=8'h10;
	15'h2aa9: q<=8'h10;
	15'h2aaa: q<=8'h48;
	15'h2aab: q<=8'h48;
	15'h2aac: q<=8'h94;
	15'h2aad: q<=8'hb0;
	15'h2aae: q<=8'hb8;
	15'h2aaf: q<=8'ha7;
	15'h2ab0: q<=8'ha7;
	15'h2ab1: q<=8'hb8;
	15'h2ab2: q<=8'hb0;
	15'h2ab3: q<=8'h94;
	15'h2ab4: q<=8'h6c;
	15'h2ab5: q<=8'h50;
	15'h2ab6: q<=8'h48;
	15'h2ab7: q<=8'h59;
	15'h2ab8: q<=8'h59;
	15'h2ab9: q<=8'h48;
	15'h2aba: q<=8'h50;
	15'h2abb: q<=8'h6c;
	15'h2abc: q<=8'h96;
	15'h2abd: q<=8'ha3;
	15'h2abe: q<=8'hc5;
	15'h2abf: q<=8'hf0;
	15'h2ac0: q<=8'hf0;
	15'h2ac1: q<=8'hc5;
	15'h2ac2: q<=8'ha3;
	15'h2ac3: q<=8'h96;
	15'h2ac4: q<=8'h6a;
	15'h2ac5: q<=8'h5d;
	15'h2ac6: q<=8'h3b;
	15'h2ac7: q<=8'h10;
	15'h2ac8: q<=8'h10;
	15'h2ac9: q<=8'h3b;
	15'h2aca: q<=8'h5d;
	15'h2acb: q<=8'h6a;
	15'h2acc: q<=8'h3d;
	15'h2acd: q<=8'h6a;
	15'h2ace: q<=8'h97;
	15'h2acf: q<=8'hc4;
	15'h2ad0: q<=8'hf0;
	15'h2ad1: q<=8'hc4;
	15'h2ad2: q<=8'h97;
	15'h2ad3: q<=8'h6a;
	15'h2ad4: q<=8'h3d;
	15'h2ad5: q<=8'h10;
	15'h2ad6: q<=8'h10;
	15'h2ad7: q<=8'h10;
	15'h2ad8: q<=8'h10;
	15'h2ad9: q<=8'h10;
	15'h2ada: q<=8'h10;
	15'h2adb: q<=8'h10;
	15'h2adc: q<=8'ha0;
	15'h2add: q<=8'he0;
	15'h2ade: q<=8'hea;
	15'h2adf: q<=8'hb0;
	15'h2ae0: q<=8'hea;
	15'h2ae1: q<=8'he0;
	15'h2ae2: q<=8'ha0;
	15'h2ae3: q<=8'h80;
	15'h2ae4: q<=8'h60;
	15'h2ae5: q<=8'h20;
	15'h2ae6: q<=8'h16;
	15'h2ae7: q<=8'h50;
	15'h2ae8: q<=8'h16;
	15'h2ae9: q<=8'h20;
	15'h2aea: q<=8'h60;
	15'h2aeb: q<=8'h80;
	15'h2aec: q<=8'hf0;
	15'h2aed: q<=8'hd0;
	15'h2aee: q<=8'hb0;
	15'h2aef: q<=8'h90;
	15'h2af0: q<=8'h70;
	15'h2af1: q<=8'h50;
	15'h2af2: q<=8'h30;
	15'h2af3: q<=8'h10;
	15'h2af4: q<=8'h10;
	15'h2af5: q<=8'h30;
	15'h2af6: q<=8'h50;
	15'h2af7: q<=8'h70;
	15'h2af8: q<=8'h90;
	15'h2af9: q<=8'hb0;
	15'h2afa: q<=8'hd0;
	15'h2afb: q<=8'hf0;
	15'h2afc: q<=8'h40;
	15'h2afd: q<=8'h40;
	15'h2afe: q<=8'h40;
	15'h2aff: q<=8'h40;
	15'h2b00: q<=8'h40;
	15'h2b01: q<=8'h40;
	15'h2b02: q<=8'h40;
	15'h2b03: q<=8'h40;
	15'h2b04: q<=8'h40;
	15'h2b05: q<=8'h40;
	15'h2b06: q<=8'h40;
	15'h2b07: q<=8'h40;
	15'h2b08: q<=8'h40;
	15'h2b09: q<=8'h40;
	15'h2b0a: q<=8'h40;
	15'h2b0b: q<=8'h40;
	15'h2b0c: q<=8'hf0;
	15'h2b0d: q<=8'hcb;
	15'h2b0e: q<=8'ha6;
	15'h2b0f: q<=8'h80;
	15'h2b10: q<=8'h5c;
	15'h2b11: q<=8'h39;
	15'h2b12: q<=8'h20;
	15'h2b13: q<=8'h12;
	15'h2b14: q<=8'h12;
	15'h2b15: q<=8'h20;
	15'h2b16: q<=8'h39;
	15'h2b17: q<=8'h5c;
	15'h2b18: q<=8'h80;
	15'h2b19: q<=8'ha6;
	15'h2b1a: q<=8'hcb;
	15'h2b1b: q<=8'hf0;
	15'h2b1c: q<=8'hc0;
	15'h2b1d: q<=8'ha6;
	15'h2b1e: q<=8'h8a;
	15'h2b1f: q<=8'h6a;
	15'h2b20: q<=8'h4a;
	15'h2b21: q<=8'h2f;
	15'h2b22: q<=8'h14;
	15'h2b23: q<=8'h24;
	15'h2b24: q<=8'h20;
	15'h2b25: q<=8'h39;
	15'h2b26: q<=8'h59;
	15'h2b27: q<=8'h75;
	15'h2b28: q<=8'h72;
	15'h2b29: q<=8'h90;
	15'h2b2a: q<=8'hb0;
	15'h2b2b: q<=8'hd0;
	15'h2b2c: q<=8'h80;
	15'h2b2d: q<=8'h57;
	15'h2b2e: q<=8'h48;
	15'h2b2f: q<=8'h57;
	15'h2b30: q<=8'h80;
	15'h2b31: q<=8'ha9;
	15'h2b32: q<=8'hba;
	15'h2b33: q<=8'ha9;
	15'h2b34: q<=8'h80;
	15'h2b35: q<=8'h57;
	15'h2b36: q<=8'h48;
	15'h2b37: q<=8'h57;
	15'h2b38: q<=8'h80;
	15'h2b39: q<=8'ha9;
	15'h2b3a: q<=8'hba;
	15'h2b3b: q<=8'ha9;
	15'h2b3c: q<=8'he4;
	15'h2b3d: q<=8'he8;
	15'h2b3e: q<=8'hb7;
	15'h2b3f: q<=8'h80;
	15'h2b40: q<=8'hb7;
	15'h2b41: q<=8'he8;
	15'h2b42: q<=8'he4;
	15'h2b43: q<=8'hb2;
	15'h2b44: q<=8'h7a;
	15'h2b45: q<=8'h47;
	15'h2b46: q<=8'h20;
	15'h2b47: q<=8'h10;
	15'h2b48: q<=8'h20;
	15'h2b49: q<=8'h47;
	15'h2b4a: q<=8'h7a;
	15'h2b4b: q<=8'hb2;
	15'h2b4c: q<=8'h90;
	15'h2b4d: q<=8'h70;
	15'h2b4e: q<=8'h70;
	15'h2b4f: q<=8'h50;
	15'h2b50: q<=8'h50;
	15'h2b51: q<=8'h30;
	15'h2b52: q<=8'h30;
	15'h2b53: q<=8'h10;
	15'h2b54: q<=8'h10;
	15'h2b55: q<=8'h30;
	15'h2b56: q<=8'h30;
	15'h2b57: q<=8'h50;
	15'h2b58: q<=8'h50;
	15'h2b59: q<=8'h70;
	15'h2b5a: q<=8'h70;
	15'h2b5b: q<=8'h90;
	15'h2b5c: q<=8'he6;
	15'h2b5d: q<=8'hd0;
	15'h2b5e: q<=8'he6;
	15'h2b5f: q<=8'hb9;
	15'h2b60: q<=8'hae;
	15'h2b61: q<=8'h80;
	15'h2b62: q<=8'h52;
	15'h2b63: q<=8'h47;
	15'h2b64: q<=8'h14;
	15'h2b65: q<=8'h30;
	15'h2b66: q<=8'h14;
	15'h2b67: q<=8'h47;
	15'h2b68: q<=8'h52;
	15'h2b69: q<=8'h80;
	15'h2b6a: q<=8'hae;
	15'h2b6b: q<=8'hb9;
	15'h2b6c: q<=8'h7e;
	15'h2b6d: q<=8'h6a;
	15'h2b6e: q<=8'h51;
	15'h2b6f: q<=8'h3a;
	15'h2b70: q<=8'h2c;
	15'h2b71: q<=8'h2c;
	15'h2b72: q<=8'h38;
	15'h2b73: q<=8'h4e;
	15'h2b74: q<=8'h4e;
	15'h2b75: q<=8'h38;
	15'h2b76: q<=8'h2c;
	15'h2b77: q<=8'h2c;
	15'h2b78: q<=8'h3a;
	15'h2b79: q<=8'h51;
	15'h2b7a: q<=8'h6a;
	15'h2b7b: q<=8'h7e;
	15'h2b7c: q<=8'h05;
	15'h2b7d: q<=8'h06;
	15'h2b7e: q<=8'h07;
	15'h2b7f: q<=8'h08;
	15'h2b80: q<=8'h09;
	15'h2b81: q<=8'h0a;
	15'h2b82: q<=8'h0b;
	15'h2b83: q<=8'h0c;
	15'h2b84: q<=8'h0d;
	15'h2b85: q<=8'h0e;
	15'h2b86: q<=8'h0f;
	15'h2b87: q<=8'h00;
	15'h2b88: q<=8'h01;
	15'h2b89: q<=8'h02;
	15'h2b8a: q<=8'h03;
	15'h2b8b: q<=8'h04;
	15'h2b8c: q<=8'h04;
	15'h2b8d: q<=8'h04;
	15'h2b8e: q<=8'h08;
	15'h2b8f: q<=8'h08;
	15'h2b90: q<=8'h08;
	15'h2b91: q<=8'h08;
	15'h2b92: q<=8'h0c;
	15'h2b93: q<=8'h0c;
	15'h2b94: q<=8'h0c;
	15'h2b95: q<=8'h0c;
	15'h2b96: q<=8'h00;
	15'h2b97: q<=8'h00;
	15'h2b98: q<=8'h00;
	15'h2b99: q<=8'h00;
	15'h2b9a: q<=8'h04;
	15'h2b9b: q<=8'h04;
	15'h2b9c: q<=8'h04;
	15'h2b9d: q<=8'h08;
	15'h2b9e: q<=8'h04;
	15'h2b9f: q<=8'h08;
	15'h2ba0: q<=8'h08;
	15'h2ba1: q<=8'h0c;
	15'h2ba2: q<=8'h08;
	15'h2ba3: q<=8'h0c;
	15'h2ba4: q<=8'h0c;
	15'h2ba5: q<=8'h00;
	15'h2ba6: q<=8'h0c;
	15'h2ba7: q<=8'h00;
	15'h2ba8: q<=8'h00;
	15'h2ba9: q<=8'h04;
	15'h2baa: q<=8'h00;
	15'h2bab: q<=8'h04;
	15'h2bac: q<=8'h06;
	15'h2bad: q<=8'h07;
	15'h2bae: q<=8'h09;
	15'h2baf: q<=8'h08;
	15'h2bb0: q<=8'h07;
	15'h2bb1: q<=8'h09;
	15'h2bb2: q<=8'h0a;
	15'h2bb3: q<=8'h0c;
	15'h2bb4: q<=8'h0e;
	15'h2bb5: q<=8'h0f;
	15'h2bb6: q<=8'h01;
	15'h2bb7: q<=8'h00;
	15'h2bb8: q<=8'h0f;
	15'h2bb9: q<=8'h01;
	15'h2bba: q<=8'h02;
	15'h2bbb: q<=8'h04;
	15'h2bbc: q<=8'h07;
	15'h2bbd: q<=8'h06;
	15'h2bbe: q<=8'h05;
	15'h2bbf: q<=8'h08;
	15'h2bc0: q<=8'h0b;
	15'h2bc1: q<=8'h0a;
	15'h2bc2: q<=8'h09;
	15'h2bc3: q<=8'h0c;
	15'h2bc4: q<=8'h0f;
	15'h2bc5: q<=8'h0e;
	15'h2bc6: q<=8'h0d;
	15'h2bc7: q<=8'h00;
	15'h2bc8: q<=8'h03;
	15'h2bc9: q<=8'h02;
	15'h2bca: q<=8'h01;
	15'h2bcb: q<=8'h04;
	15'h2bcc: q<=8'h05;
	15'h2bcd: q<=8'h05;
	15'h2bce: q<=8'h05;
	15'h2bcf: q<=8'h05;
	15'h2bd0: q<=8'h0b;
	15'h2bd1: q<=8'h0b;
	15'h2bd2: q<=8'h0b;
	15'h2bd3: q<=8'h0b;
	15'h2bd4: q<=8'h0b;
	15'h2bd5: q<=8'h00;
	15'h2bd6: q<=8'h00;
	15'h2bd7: q<=8'h00;
	15'h2bd8: q<=8'h00;
	15'h2bd9: q<=8'h00;
	15'h2bda: q<=8'h00;
	15'h2bdb: q<=8'h05;
	15'h2bdc: q<=8'h04;
	15'h2bdd: q<=8'h08;
	15'h2bde: q<=8'h0b;
	15'h2bdf: q<=8'h05;
	15'h2be0: q<=8'h08;
	15'h2be1: q<=8'h0c;
	15'h2be2: q<=8'h0e;
	15'h2be3: q<=8'h09;
	15'h2be4: q<=8'h0c;
	15'h2be5: q<=8'h00;
	15'h2be6: q<=8'h03;
	15'h2be7: q<=8'h0d;
	15'h2be8: q<=8'h00;
	15'h2be9: q<=8'h04;
	15'h2bea: q<=8'h07;
	15'h2beb: q<=8'h02;
	15'h2bec: q<=8'h0d;
	15'h2bed: q<=8'h0d;
	15'h2bee: q<=8'h0d;
	15'h2bef: q<=8'h0d;
	15'h2bf0: q<=8'h0d;
	15'h2bf1: q<=8'h0d;
	15'h2bf2: q<=8'h0d;
	15'h2bf3: q<=8'h00;
	15'h2bf4: q<=8'h03;
	15'h2bf5: q<=8'h03;
	15'h2bf6: q<=8'h03;
	15'h2bf7: q<=8'h03;
	15'h2bf8: q<=8'h03;
	15'h2bf9: q<=8'h03;
	15'h2bfa: q<=8'h03;
	15'h2bfb: q<=8'h00;
	15'h2bfc: q<=8'h00;
	15'h2bfd: q<=8'h00;
	15'h2bfe: q<=8'h00;
	15'h2bff: q<=8'h00;
	15'h2c00: q<=8'h00;
	15'h2c01: q<=8'h00;
	15'h2c02: q<=8'h00;
	15'h2c03: q<=8'h00;
	15'h2c04: q<=8'h00;
	15'h2c05: q<=8'h00;
	15'h2c06: q<=8'h00;
	15'h2c07: q<=8'h00;
	15'h2c08: q<=8'h00;
	15'h2c09: q<=8'h00;
	15'h2c0a: q<=8'h00;
	15'h2c0b: q<=8'h00;
	15'h2c0c: q<=8'h0c;
	15'h2c0d: q<=8'h0c;
	15'h2c0e: q<=8'h0c;
	15'h2c0f: q<=8'h0d;
	15'h2c10: q<=8'h0e;
	15'h2c11: q<=8'h0f;
	15'h2c12: q<=8'h0f;
	15'h2c13: q<=8'h00;
	15'h2c14: q<=8'h01;
	15'h2c15: q<=8'h01;
	15'h2c16: q<=8'h02;
	15'h2c17: q<=8'h03;
	15'h2c18: q<=8'h04;
	15'h2c19: q<=8'h04;
	15'h2c1a: q<=8'h04;
	15'h2c1b: q<=8'h00;
	15'h2c1c: q<=8'h0e;
	15'h2c1d: q<=8'h0d;
	15'h2c1e: q<=8'h0c;
	15'h2c1f: q<=8'h0d;
	15'h2c20: q<=8'h0d;
	15'h2c21: q<=8'h0d;
	15'h2c22: q<=8'h01;
	15'h2c23: q<=8'h0f;
	15'h2c24: q<=8'h02;
	15'h2c25: q<=8'h03;
	15'h2c26: q<=8'h03;
	15'h2c27: q<=8'h00;
	15'h2c28: q<=8'h03;
	15'h2c29: q<=8'h03;
	15'h2c2a: q<=8'h03;
	15'h2c2b: q<=8'h00;
	15'h2c2c: q<=8'h0b;
	15'h2c2d: q<=8'h09;
	15'h2c2e: q<=8'h07;
	15'h2c2f: q<=8'h05;
	15'h2c30: q<=8'h03;
	15'h2c31: q<=8'h01;
	15'h2c32: q<=8'h0f;
	15'h2c33: q<=8'h0d;
	15'h2c34: q<=8'h0d;
	15'h2c35: q<=8'h0f;
	15'h2c36: q<=8'h01;
	15'h2c37: q<=8'h03;
	15'h2c38: q<=8'h05;
	15'h2c39: q<=8'h07;
	15'h2c3a: q<=8'h09;
	15'h2c3b: q<=8'h0b;
	15'h2c3c: q<=8'h08;
	15'h2c3d: q<=8'h0b;
	15'h2c3e: q<=8'h0c;
	15'h2c3f: q<=8'h04;
	15'h2c40: q<=8'h05;
	15'h2c41: q<=8'h08;
	15'h2c42: q<=8'h0b;
	15'h2c43: q<=8'h0c;
	15'h2c44: q<=8'h0d;
	15'h2c45: q<=8'h0e;
	15'h2c46: q<=8'h0f;
	15'h2c47: q<=8'h01;
	15'h2c48: q<=8'h02;
	15'h2c49: q<=8'h03;
	15'h2c4a: q<=8'h04;
	15'h2c4b: q<=8'h05;
	15'h2c4c: q<=8'h0c;
	15'h2c4d: q<=8'h00;
	15'h2c4e: q<=8'h0c;
	15'h2c4f: q<=8'h00;
	15'h2c50: q<=8'h0c;
	15'h2c51: q<=8'h00;
	15'h2c52: q<=8'h0c;
	15'h2c53: q<=8'h00;
	15'h2c54: q<=8'h04;
	15'h2c55: q<=8'h00;
	15'h2c56: q<=8'h04;
	15'h2c57: q<=8'h00;
	15'h2c58: q<=8'h04;
	15'h2c59: q<=8'h00;
	15'h2c5a: q<=8'h04;
	15'h2c5b: q<=8'h00;
	15'h2c5c: q<=8'h0a;
	15'h2c5d: q<=8'h06;
	15'h2c5e: q<=8'h0c;
	15'h2c5f: q<=8'h08;
	15'h2c60: q<=8'h0e;
	15'h2c61: q<=8'h0a;
	15'h2c62: q<=8'h00;
	15'h2c63: q<=8'h0c;
	15'h2c64: q<=8'h02;
	15'h2c65: q<=8'h0e;
	15'h2c66: q<=8'h04;
	15'h2c67: q<=8'h00;
	15'h2c68: q<=8'h06;
	15'h2c69: q<=8'h02;
	15'h2c6a: q<=8'h08;
	15'h2c6b: q<=8'h04;
	15'h2c6c: q<=8'h0e;
	15'h2c6d: q<=8'h0c;
	15'h2c6e: q<=8'h0d;
	15'h2c6f: q<=8'h0e;
	15'h2c70: q<=8'h00;
	15'h2c71: q<=8'h02;
	15'h2c72: q<=8'h02;
	15'h2c73: q<=8'h00;
	15'h2c74: q<=8'h0e;
	15'h2c75: q<=8'h0e;
	15'h2c76: q<=8'h00;
	15'h2c77: q<=8'h02;
	15'h2c78: q<=8'h03;
	15'h2c79: q<=8'h04;
	15'h2c7a: q<=8'h02;
	15'h2c7b: q<=8'h00;
	15'h2c7c: q<=8'h00;
	15'h2c7d: q<=8'h01;
	15'h2c7e: q<=8'h02;
	15'h2c7f: q<=8'h03;
	15'h2c80: q<=8'h04;
	15'h2c81: q<=8'h05;
	15'h2c82: q<=8'h06;
	15'h2c83: q<=8'h07;
	15'h2c84: q<=8'h0d;
	15'h2c85: q<=8'h09;
	15'h2c86: q<=8'h08;
	15'h2c87: q<=8'h0c;
	15'h2c88: q<=8'h0e;
	15'h2c89: q<=8'h0f;
	15'h2c8a: q<=8'h0a;
	15'h2c8b: q<=8'h0b;
	15'h2c8c: q<=8'h18;
	15'h2c8d: q<=8'h1c;
	15'h2c8e: q<=8'h18;
	15'h2c8f: q<=8'h0f;
	15'h2c90: q<=8'h18;
	15'h2c91: q<=8'h18;
	15'h2c92: q<=8'h18;
	15'h2c93: q<=8'h18;
	15'h2c94: q<=8'h0a;
	15'h2c95: q<=8'h18;
	15'h2c96: q<=8'h10;
	15'h2c97: q<=8'h0f;
	15'h2c98: q<=8'h18;
	15'h2c99: q<=8'h0c;
	15'h2c9a: q<=8'h14;
	15'h2c9b: q<=8'h0a;
	15'h2c9c: q<=8'h50;
	15'h2c9d: q<=8'h50;
	15'h2c9e: q<=8'h50;
	15'h2c9f: q<=8'h68;
	15'h2ca0: q<=8'h50;
	15'h2ca1: q<=8'h50;
	15'h2ca2: q<=8'h68;
	15'h2ca3: q<=8'hb0;
	15'h2ca4: q<=8'ha0;
	15'h2ca5: q<=8'h50;
	15'h2ca6: q<=8'h90;
	15'h2ca7: q<=8'h80;
	15'h2ca8: q<=8'h20;
	15'h2ca9: q<=8'hb0;
	15'h2caa: q<=8'h60;
	15'h2cab: q<=8'ha0;
	15'h2cac: q<=8'h40;
	15'h2cad: q<=8'h20;
	15'h2cae: q<=8'h40;
	15'h2caf: q<=8'h80;
	15'h2cb0: q<=8'h40;
	15'h2cb1: q<=8'h40;
	15'h2cb2: q<=8'h70;
	15'h2cb3: q<=8'h60;
	15'h2cb4: q<=8'h00;
	15'h2cb5: q<=8'h20;
	15'h2cb6: q<=8'h40;
	15'h2cb7: q<=8'h00;
	15'h2cb8: q<=8'ha0;
	15'h2cb9: q<=8'h40;
	15'h2cba: q<=8'h40;
	15'h2cbb: q<=8'h00;
	15'h2cbc: q<=8'hff;
	15'h2cbd: q<=8'hff;
	15'h2cbe: q<=8'hff;
	15'h2cbf: q<=8'hff;
	15'h2cc0: q<=8'hff;
	15'h2cc1: q<=8'hff;
	15'h2cc2: q<=8'hff;
	15'h2cc3: q<=8'h00;
	15'h2cc4: q<=8'h01;
	15'h2cc5: q<=8'hff;
	15'h2cc6: q<=8'h00;
	15'h2cc7: q<=8'h00;
	15'h2cc8: q<=8'hfe;
	15'h2cc9: q<=8'h01;
	15'h2cca: q<=8'hff;
	15'h2ccb: q<=8'h01;
	15'h2ccc: q<=8'h00;
	15'h2ccd: q<=8'h00;
	15'h2cce: q<=8'h00;
	15'h2ccf: q<=8'h00;
	15'h2cd0: q<=8'h00;
	15'h2cd1: q<=8'h00;
	15'h2cd2: q<=8'h00;
	15'h2cd3: q<=8'hff;
	15'h2cd4: q<=8'hff;
	15'h2cd5: q<=8'hff;
	15'h2cd6: q<=8'hff;
	15'h2cd7: q<=8'h00;
	15'h2cd8: q<=8'h00;
	15'h2cd9: q<=8'hff;
	15'h2cda: q<=8'h00;
	15'h2cdb: q<=8'hff;
	15'h2cdc: q<=8'h00;
	15'h2cdd: q<=8'h00;
	15'h2cde: q<=8'h60;
	15'h2cdf: q<=8'h40;
	15'h2ce0: q<=8'h00;
	15'h2ce1: q<=8'h00;
	15'h2ce2: q<=8'h48;
	15'h2ce3: q<=8'h40;
	15'h2ce4: q<=8'h50;
	15'h2ce5: q<=8'h28;
	15'h2ce6: q<=8'h50;
	15'h2ce7: q<=8'h00;
	15'h2ce8: q<=8'h00;
	15'h2ce9: q<=8'h50;
	15'h2cea: q<=8'h00;
	15'h2ceb: q<=8'h40;
	15'h2cec: q<=8'h04;
	15'h2ced: q<=8'h04;
	15'h2cee: q<=8'h03;
	15'h2cef: q<=8'h04;
	15'h2cf0: q<=8'h04;
	15'h2cf1: q<=8'h04;
	15'h2cf2: q<=8'h03;
	15'h2cf3: q<=8'h04;
	15'h2cf4: q<=8'h05;
	15'h2cf5: q<=8'h04;
	15'h2cf6: q<=8'h04;
	15'h2cf7: q<=8'h04;
	15'h2cf8: q<=8'h04;
	15'h2cf9: q<=8'h04;
	15'h2cfa: q<=8'h04;
	15'h2cfb: q<=8'h05;
	15'h2cfc: q<=8'h3e;
	15'h2cfd: q<=8'h85;
	15'h2cfe: q<=8'h55;
	15'h2cff: q<=8'hb9;
	15'h2d00: q<=8'h35;
	15'h2d01: q<=8'h04;
	15'h2d02: q<=8'h85;
	15'h2d03: q<=8'h56;
	15'h2d04: q<=8'hb9;
	15'h2d05: q<=8'h45;
	15'h2d06: q<=8'h04;
	15'h2d07: q<=8'h85;
	15'h2d08: q<=8'h58;
	15'h2d09: q<=8'h20;
	15'h2d0a: q<=8'h98;
	15'h2d0b: q<=8'hc0;
	15'h2d0c: q<=8'ha2;
	15'h2d0d: q<=8'h61;
	15'h2d0e: q<=8'h20;
	15'h2d0f: q<=8'h65;
	15'h2d10: q<=8'hc7;
	15'h2d11: q<=8'ha9;
	15'h2d12: q<=8'h00;
	15'h2d13: q<=8'h85;
	15'h2d14: q<=8'ha9;
	15'h2d15: q<=8'h20;
	15'h2d16: q<=8'h3e;
	15'h2d17: q<=8'hbd;
	15'h2d18: q<=8'ha5;
	15'h2d19: q<=8'h78;
	15'h2d1a: q<=8'h49;
	15'h2d1b: q<=8'h07;
	15'h2d1c: q<=8'h0a;
	15'h2d1d: q<=8'hc9;
	15'h2d1e: q<=8'h0a;
	15'h2d1f: q<=8'hb0;
	15'h2d20: q<=8'h02;
	15'h2d21: q<=8'ha9;
	15'h2d22: q<=8'h0a;
	15'h2d23: q<=8'h0a;
	15'h2d24: q<=8'h0a;
	15'h2d25: q<=8'h0a;
	15'h2d26: q<=8'h0a;
	15'h2d27: q<=8'h91;
	15'h2d28: q<=8'h74;
	15'h2d29: q<=8'hc8;
	15'h2d2a: q<=8'ha9;
	15'h2d2b: q<=8'h60;
	15'h2d2c: q<=8'h91;
	15'h2d2d: q<=8'h74;
	15'h2d2e: q<=8'hc8;
	15'h2d2f: q<=8'h84;
	15'h2d30: q<=8'ha9;
	15'h2d31: q<=8'ha4;
	15'h2d32: q<=8'h55;
	15'h2d33: q<=8'hbe;
	15'h2d34: q<=8'hc9;
	15'h2d35: q<=8'hce;
	15'h2d36: q<=8'hb9;
	15'h2d37: q<=8'hc8;
	15'h2d38: q<=8'hce;
	15'h2d39: q<=8'ha4;
	15'h2d3a: q<=8'ha9;
	15'h2d3b: q<=8'h4c;
	15'h2d3c: q<=8'h59;
	15'h2d3d: q<=8'hdf;
	15'h2d3e: q<=8'ha5;
	15'h2d3f: q<=8'h57;
	15'h2d40: q<=8'hc9;
	15'h2d41: q<=8'h10;
	15'h2d42: q<=8'h90;
	15'h2d43: q<=8'h48;
	15'h2d44: q<=8'h38;
	15'h2d45: q<=8'he5;
	15'h2d46: q<=8'h5f;
	15'h2d47: q<=8'h8d;
	15'h2d48: q<=8'h95;
	15'h2d49: q<=8'h60;
	15'h2d4a: q<=8'ha9;
	15'h2d4b: q<=8'h00;
	15'h2d4c: q<=8'he5;
	15'h2d4d: q<=8'h5b;
	15'h2d4e: q<=8'h8d;
	15'h2d4f: q<=8'h96;
	15'h2d50: q<=8'h60;
	15'h2d51: q<=8'ha9;
	15'h2d52: q<=8'h18;
	15'h2d53: q<=8'h8d;
	15'h2d54: q<=8'h8c;
	15'h2d55: q<=8'h60;
	15'h2d56: q<=8'ha5;
	15'h2d57: q<=8'ha0;
	15'h2d58: q<=8'h8d;
	15'h2d59: q<=8'h8e;
	15'h2d5a: q<=8'h60;
	15'h2d5b: q<=8'h8d;
	15'h2d5c: q<=8'h94;
	15'h2d5d: q<=8'h60;
	15'h2d5e: q<=8'h2c;
	15'h2d5f: q<=8'h40;
	15'h2d60: q<=8'h60;
	15'h2d61: q<=8'h30;
	15'h2d62: q<=8'hfb;
	15'h2d63: q<=8'had;
	15'h2d64: q<=8'h60;
	15'h2d65: q<=8'h60;
	15'h2d66: q<=8'h85;
	15'h2d67: q<=8'h79;
	15'h2d68: q<=8'had;
	15'h2d69: q<=8'h70;
	15'h2d6a: q<=8'h60;
	15'h2d6b: q<=8'h85;
	15'h2d6c: q<=8'h7a;
	15'h2d6d: q<=8'ha2;
	15'h2d6e: q<=8'h0f;
	15'h2d6f: q<=8'h8e;
	15'h2d70: q<=8'h8c;
	15'h2d71: q<=8'h60;
	15'h2d72: q<=8'h38;
	15'h2d73: q<=8'he9;
	15'h2d74: q<=8'h01;
	15'h2d75: q<=8'hd0;
	15'h2d76: q<=8'h02;
	15'h2d77: q<=8'ha9;
	15'h2d78: q<=8'h01;
	15'h2d79: q<=8'ha2;
	15'h2d7a: q<=8'h00;
	15'h2d7b: q<=8'he8;
	15'h2d7c: q<=8'h06;
	15'h2d7d: q<=8'h79;
	15'h2d7e: q<=8'h2a;
	15'h2d7f: q<=8'h90;
	15'h2d80: q<=8'hfa;
	15'h2d81: q<=8'h4a;
	15'h2d82: q<=8'h49;
	15'h2d83: q<=8'h7f;
	15'h2d84: q<=8'h18;
	15'h2d85: q<=8'h69;
	15'h2d86: q<=8'h01;
	15'h2d87: q<=8'ha8;
	15'h2d88: q<=8'h8a;
	15'h2d89: q<=8'hb8;
	15'h2d8a: q<=8'h50;
	15'h2d8b: q<=8'h04;
	15'h2d8c: q<=8'ha9;
	15'h2d8d: q<=8'h01;
	15'h2d8e: q<=8'ha0;
	15'h2d8f: q<=8'h00;
	15'h2d90: q<=8'h85;
	15'h2d91: q<=8'h78;
	15'h2d92: q<=8'h48;
	15'h2d93: q<=8'h98;
	15'h2d94: q<=8'ha4;
	15'h2d95: q<=8'ha9;
	15'h2d96: q<=8'h91;
	15'h2d97: q<=8'h74;
	15'h2d98: q<=8'hc8;
	15'h2d99: q<=8'h68;
	15'h2d9a: q<=8'h09;
	15'h2d9b: q<=8'h70;
	15'h2d9c: q<=8'h91;
	15'h2d9d: q<=8'h74;
	15'h2d9e: q<=8'hc8;
	15'h2d9f: q<=8'h60;
	15'h2da0: q<=8'h85;
	15'h2da1: q<=8'h36;
	15'h2da2: q<=8'hb9;
	15'h2da3: q<=8'hce;
	15'h2da4: q<=8'h03;
	15'h2da5: q<=8'h85;
	15'h2da6: q<=8'h56;
	15'h2da7: q<=8'hb9;
	15'h2da8: q<=8'hde;
	15'h2da9: q<=8'h03;
	15'h2daa: q<=8'h85;
	15'h2dab: q<=8'h58;
	15'h2dac: q<=8'ha5;
	15'h2dad: q<=8'h57;
	15'h2dae: q<=8'h85;
	15'h2daf: q<=8'h2f;
	15'h2db0: q<=8'h98;
	15'h2db1: q<=8'h18;
	15'h2db2: q<=8'h69;
	15'h2db3: q<=8'h01;
	15'h2db4: q<=8'h29;
	15'h2db5: q<=8'h0f;
	15'h2db6: q<=8'haa;
	15'h2db7: q<=8'hbd;
	15'h2db8: q<=8'hce;
	15'h2db9: q<=8'h03;
	15'h2dba: q<=8'h85;
	15'h2dbb: q<=8'h2e;
	15'h2dbc: q<=8'hbd;
	15'h2dbd: q<=8'hde;
	15'h2dbe: q<=8'h03;
	15'h2dbf: q<=8'h85;
	15'h2dc0: q<=8'h30;
	15'h2dc1: q<=8'ha9;
	15'h2dc2: q<=8'h00;
	15'h2dc3: q<=8'h85;
	15'h2dc4: q<=8'h59;
	15'h2dc5: q<=8'ha9;
	15'h2dc6: q<=8'h04;
	15'h2dc7: q<=8'h85;
	15'h2dc8: q<=8'h5a;
	15'h2dc9: q<=8'ha4;
	15'h2dca: q<=8'h36;
	15'h2dcb: q<=8'ha5;
	15'h2dcc: q<=8'h5b;
	15'h2dcd: q<=8'h30;
	15'h2dce: q<=8'h07;
	15'h2dcf: q<=8'ha5;
	15'h2dd0: q<=8'h57;
	15'h2dd1: q<=8'hc5;
	15'h2dd2: q<=8'h5f;
	15'h2dd3: q<=8'hb0;
	15'h2dd4: q<=8'h01;
	15'h2dd5: q<=8'h60;
	15'h2dd6: q<=8'hb9;
	15'h2dd7: q<=8'hb6;
	15'h2dd8: q<=8'hbf;
	15'h2dd9: q<=8'h85;
	15'h2dda: q<=8'h99;
	15'h2ddb: q<=8'hb9;
	15'h2ddc: q<=8'hc4;
	15'h2ddd: q<=8'hbf;
	15'h2dde: q<=8'h85;
	15'h2ddf: q<=8'h38;
	15'h2de0: q<=8'ha4;
	15'h2de1: q<=8'h9e;
	15'h2de2: q<=8'ha9;
	15'h2de3: q<=8'h08;
	15'h2de4: q<=8'h20;
	15'h2de5: q<=8'h4c;
	15'h2de6: q<=8'hdf;
	15'h2de7: q<=8'h20;
	15'h2de8: q<=8'h98;
	15'h2de9: q<=8'hc0;
	15'h2dea: q<=8'ha2;
	15'h2deb: q<=8'h61;
	15'h2dec: q<=8'h20;
	15'h2ded: q<=8'h65;
	15'h2dee: q<=8'hc7;
	15'h2def: q<=8'ha5;
	15'h2df0: q<=8'h2e;
	15'h2df1: q<=8'h85;
	15'h2df2: q<=8'h56;
	15'h2df3: q<=8'ha5;
	15'h2df4: q<=8'h2f;
	15'h2df5: q<=8'h85;
	15'h2df6: q<=8'h57;
	15'h2df7: q<=8'ha5;
	15'h2df8: q<=8'h30;
	15'h2df9: q<=8'h85;
	15'h2dfa: q<=8'h58;
	15'h2dfb: q<=8'h20;
	15'h2dfc: q<=8'h98;
	15'h2dfd: q<=8'hc0;
	15'h2dfe: q<=8'ha4;
	15'h2dff: q<=8'h59;
	15'h2e00: q<=8'ha5;
	15'h2e01: q<=8'h5a;
	15'h2e02: q<=8'h20;
	15'h2e03: q<=8'h6c;
	15'h2e04: q<=8'hdf;
	15'h2e05: q<=8'ha5;
	15'h2e06: q<=8'h61;
	15'h2e07: q<=8'h38;
	15'h2e08: q<=8'he5;
	15'h2e09: q<=8'h6a;
	15'h2e0a: q<=8'h85;
	15'h2e0b: q<=8'h79;
	15'h2e0c: q<=8'ha5;
	15'h2e0d: q<=8'h62;
	15'h2e0e: q<=8'he5;
	15'h2e0f: q<=8'h6b;
	15'h2e10: q<=8'h85;
	15'h2e11: q<=8'h9b;
	15'h2e12: q<=8'h30;
	15'h2e13: q<=8'h09;
	15'h2e14: q<=8'hf0;
	15'h2e15: q<=8'h04;
	15'h2e16: q<=8'ha9;
	15'h2e17: q<=8'hff;
	15'h2e18: q<=8'h85;
	15'h2e19: q<=8'h79;
	15'h2e1a: q<=8'hb8;
	15'h2e1b: q<=8'h50;
	15'h2e1c: q<=8'h16;
	15'h2e1d: q<=8'hc9;
	15'h2e1e: q<=8'hff;
	15'h2e1f: q<=8'hf0;
	15'h2e20: q<=8'h05;
	15'h2e21: q<=8'ha9;
	15'h2e22: q<=8'hff;
	15'h2e23: q<=8'hb8;
	15'h2e24: q<=8'h50;
	15'h2e25: q<=8'h0b;
	15'h2e26: q<=8'ha5;
	15'h2e27: q<=8'h79;
	15'h2e28: q<=8'h49;
	15'h2e29: q<=8'hff;
	15'h2e2a: q<=8'h18;
	15'h2e2b: q<=8'h69;
	15'h2e2c: q<=8'h01;
	15'h2e2d: q<=8'h90;
	15'h2e2e: q<=8'h02;
	15'h2e2f: q<=8'ha9;
	15'h2e30: q<=8'hff;
	15'h2e31: q<=8'h85;
	15'h2e32: q<=8'h79;
	15'h2e33: q<=8'ha5;
	15'h2e34: q<=8'h63;
	15'h2e35: q<=8'h38;
	15'h2e36: q<=8'he5;
	15'h2e37: q<=8'h6c;
	15'h2e38: q<=8'h85;
	15'h2e39: q<=8'h89;
	15'h2e3a: q<=8'ha5;
	15'h2e3b: q<=8'h64;
	15'h2e3c: q<=8'he5;
	15'h2e3d: q<=8'h6d;
	15'h2e3e: q<=8'h85;
	15'h2e3f: q<=8'h9d;
	15'h2e40: q<=8'h30;
	15'h2e41: q<=8'h09;
	15'h2e42: q<=8'hf0;
	15'h2e43: q<=8'h04;
	15'h2e44: q<=8'ha9;
	15'h2e45: q<=8'hff;
	15'h2e46: q<=8'h85;
	15'h2e47: q<=8'h89;
	15'h2e48: q<=8'hb8;
	15'h2e49: q<=8'h50;
	15'h2e4a: q<=8'h12;
	15'h2e4b: q<=8'hc9;
	15'h2e4c: q<=8'hff;
	15'h2e4d: q<=8'hf0;
	15'h2e4e: q<=8'h05;
	15'h2e4f: q<=8'ha9;
	15'h2e50: q<=8'hff;
	15'h2e51: q<=8'hb8;
	15'h2e52: q<=8'h50;
	15'h2e53: q<=8'h07;
	15'h2e54: q<=8'ha5;
	15'h2e55: q<=8'h89;
	15'h2e56: q<=8'h49;
	15'h2e57: q<=8'hff;
	15'h2e58: q<=8'h18;
	15'h2e59: q<=8'h69;
	15'h2e5a: q<=8'h01;
	15'h2e5b: q<=8'h85;
	15'h2e5c: q<=8'h89;
	15'h2e5d: q<=8'ha9;
	15'h2e5e: q<=8'h00;
	15'h2e5f: q<=8'h85;
	15'h2e60: q<=8'h82;
	15'h2e61: q<=8'h85;
	15'h2e62: q<=8'h92;
	15'h2e63: q<=8'ha5;
	15'h2e64: q<=8'h79;
	15'h2e65: q<=8'h0a;
	15'h2e66: q<=8'h26;
	15'h2e67: q<=8'h82;
	15'h2e68: q<=8'h85;
	15'h2e69: q<=8'h7a;
	15'h2e6a: q<=8'h0a;
	15'h2e6b: q<=8'h85;
	15'h2e6c: q<=8'h7c;
	15'h2e6d: q<=8'ha5;
	15'h2e6e: q<=8'h82;
	15'h2e6f: q<=8'h2a;
	15'h2e70: q<=8'h85;
	15'h2e71: q<=8'h84;
	15'h2e72: q<=8'ha5;
	15'h2e73: q<=8'h7c;
	15'h2e74: q<=8'h65;
	15'h2e75: q<=8'h79;
	15'h2e76: q<=8'h85;
	15'h2e77: q<=8'h7d;
	15'h2e78: q<=8'ha5;
	15'h2e79: q<=8'h84;
	15'h2e7a: q<=8'h69;
	15'h2e7b: q<=8'h00;
	15'h2e7c: q<=8'h85;
	15'h2e7d: q<=8'h85;
	15'h2e7e: q<=8'ha5;
	15'h2e7f: q<=8'h7a;
	15'h2e80: q<=8'h65;
	15'h2e81: q<=8'h79;
	15'h2e82: q<=8'h85;
	15'h2e83: q<=8'h7b;
	15'h2e84: q<=8'ha5;
	15'h2e85: q<=8'h82;
	15'h2e86: q<=8'h69;
	15'h2e87: q<=8'h00;
	15'h2e88: q<=8'h85;
	15'h2e89: q<=8'h83;
	15'h2e8a: q<=8'h85;
	15'h2e8b: q<=8'h86;
	15'h2e8c: q<=8'ha5;
	15'h2e8d: q<=8'h7b;
	15'h2e8e: q<=8'h0a;
	15'h2e8f: q<=8'h85;
	15'h2e90: q<=8'h7e;
	15'h2e91: q<=8'h26;
	15'h2e92: q<=8'h86;
	15'h2e93: q<=8'h65;
	15'h2e94: q<=8'h79;
	15'h2e95: q<=8'h85;
	15'h2e96: q<=8'h7f;
	15'h2e97: q<=8'ha5;
	15'h2e98: q<=8'h86;
	15'h2e99: q<=8'h69;
	15'h2e9a: q<=8'h00;
	15'h2e9b: q<=8'h85;
	15'h2e9c: q<=8'h87;
	15'h2e9d: q<=8'ha5;
	15'h2e9e: q<=8'h89;
	15'h2e9f: q<=8'h0a;
	15'h2ea0: q<=8'h26;
	15'h2ea1: q<=8'h92;
	15'h2ea2: q<=8'h85;
	15'h2ea3: q<=8'h8a;
	15'h2ea4: q<=8'h0a;
	15'h2ea5: q<=8'h85;
	15'h2ea6: q<=8'h8c;
	15'h2ea7: q<=8'ha5;
	15'h2ea8: q<=8'h92;
	15'h2ea9: q<=8'h2a;
	15'h2eaa: q<=8'h85;
	15'h2eab: q<=8'h94;
	15'h2eac: q<=8'ha5;
	15'h2ead: q<=8'h8c;
	15'h2eae: q<=8'h65;
	15'h2eaf: q<=8'h89;
	15'h2eb0: q<=8'h85;
	15'h2eb1: q<=8'h8d;
	15'h2eb2: q<=8'ha5;
	15'h2eb3: q<=8'h94;
	15'h2eb4: q<=8'h69;
	15'h2eb5: q<=8'h00;
	15'h2eb6: q<=8'h85;
	15'h2eb7: q<=8'h95;
	15'h2eb8: q<=8'ha5;
	15'h2eb9: q<=8'h8a;
	15'h2eba: q<=8'h65;
	15'h2ebb: q<=8'h89;
	15'h2ebc: q<=8'h85;
	15'h2ebd: q<=8'h8b;
	15'h2ebe: q<=8'ha5;
	15'h2ebf: q<=8'h92;
	15'h2ec0: q<=8'h69;
	15'h2ec1: q<=8'h00;
	15'h2ec2: q<=8'h85;
	15'h2ec3: q<=8'h93;
	15'h2ec4: q<=8'h85;
	15'h2ec5: q<=8'h96;
	15'h2ec6: q<=8'ha5;
	15'h2ec7: q<=8'h8b;
	15'h2ec8: q<=8'h0a;
	15'h2ec9: q<=8'h85;
	15'h2eca: q<=8'h8e;
	15'h2ecb: q<=8'h26;
	15'h2ecc: q<=8'h96;
	15'h2ecd: q<=8'h65;
	15'h2ece: q<=8'h89;
	15'h2ecf: q<=8'h85;
	15'h2ed0: q<=8'h8f;
	15'h2ed1: q<=8'ha5;
	15'h2ed2: q<=8'h96;
	15'h2ed3: q<=8'h69;
	15'h2ed4: q<=8'h00;
	15'h2ed5: q<=8'h85;
	15'h2ed6: q<=8'h97;
	15'h2ed7: q<=8'ha0;
	15'h2ed8: q<=8'h00;
	15'h2ed9: q<=8'h84;
	15'h2eda: q<=8'ha9;
	15'h2edb: q<=8'ha4;
	15'h2edc: q<=8'h38;
	15'h2edd: q<=8'hb9;
	15'h2ede: q<=8'hd3;
	15'h2edf: q<=8'hbf;
	15'h2ee0: q<=8'hc9;
	15'h2ee1: q<=8'h01;
	15'h2ee2: q<=8'hd0;
	15'h2ee3: q<=8'h02;
	15'h2ee4: q<=8'ha9;
	15'h2ee5: q<=8'hc0;
	15'h2ee6: q<=8'h85;
	15'h2ee7: q<=8'h73;
	15'h2ee8: q<=8'hb9;
	15'h2ee9: q<=8'hd2;
	15'h2eea: q<=8'hbf;
	15'h2eeb: q<=8'h85;
	15'h2eec: q<=8'h2d;
	15'h2eed: q<=8'hc8;
	15'h2eee: q<=8'hc8;
	15'h2eef: q<=8'h84;
	15'h2ef0: q<=8'h38;
	15'h2ef1: q<=8'haa;
	15'h2ef2: q<=8'h29;
	15'h2ef3: q<=8'h07;
	15'h2ef4: q<=8'ha8;
	15'h2ef5: q<=8'h8a;
	15'h2ef6: q<=8'h0a;
	15'h2ef7: q<=8'h85;
	15'h2ef8: q<=8'h2b;
	15'h2ef9: q<=8'h4a;
	15'h2efa: q<=8'h4a;
	15'h2efb: q<=8'h4a;
	15'h2efc: q<=8'h4a;
	15'h2efd: q<=8'h29;
	15'h2efe: q<=8'h07;
	15'h2eff: q<=8'haa;
	15'h2f00: q<=8'ha5;
	15'h2f01: q<=8'h2b;
	15'h2f02: q<=8'h45;
	15'h2f03: q<=8'h9b;
	15'h2f04: q<=8'h30;
	15'h2f05: q<=8'h0b;
	15'h2f06: q<=8'hb9;
	15'h2f07: q<=8'h78;
	15'h2f08: q<=8'h00;
	15'h2f09: q<=8'h85;
	15'h2f0a: q<=8'h61;
	15'h2f0b: q<=8'hb9;
	15'h2f0c: q<=8'h80;
	15'h2f0d: q<=8'h00;
	15'h2f0e: q<=8'hb8;
	15'h2f0f: q<=8'h50;
	15'h2f10: q<=8'h11;
	15'h2f11: q<=8'hb9;
	15'h2f12: q<=8'h78;
	15'h2f13: q<=8'h00;
	15'h2f14: q<=8'h49;
	15'h2f15: q<=8'hff;
	15'h2f16: q<=8'h18;
	15'h2f17: q<=8'h69;
	15'h2f18: q<=8'h01;
	15'h2f19: q<=8'h85;
	15'h2f1a: q<=8'h61;
	15'h2f1b: q<=8'hb9;
	15'h2f1c: q<=8'h80;
	15'h2f1d: q<=8'h00;
	15'h2f1e: q<=8'h49;
	15'h2f1f: q<=8'hff;
	15'h2f20: q<=8'h69;
	15'h2f21: q<=8'h00;
	15'h2f22: q<=8'h85;
	15'h2f23: q<=8'h62;
	15'h2f24: q<=8'ha5;
	15'h2f25: q<=8'h2d;
	15'h2f26: q<=8'h45;
	15'h2f27: q<=8'h9d;
	15'h2f28: q<=8'h10;
	15'h2f29: q<=8'h0e;
	15'h2f2a: q<=8'hb5;
	15'h2f2b: q<=8'h88;
	15'h2f2c: q<=8'h18;
	15'h2f2d: q<=8'h65;
	15'h2f2e: q<=8'h61;
	15'h2f2f: q<=8'h85;
	15'h2f30: q<=8'h61;
	15'h2f31: q<=8'hb5;
	15'h2f32: q<=8'h90;
	15'h2f33: q<=8'h65;
	15'h2f34: q<=8'h62;
	15'h2f35: q<=8'hb8;
	15'h2f36: q<=8'h50;
	15'h2f37: q<=8'h0b;
	15'h2f38: q<=8'ha5;
	15'h2f39: q<=8'h61;
	15'h2f3a: q<=8'h38;
	15'h2f3b: q<=8'hf5;
	15'h2f3c: q<=8'h88;
	15'h2f3d: q<=8'h85;
	15'h2f3e: q<=8'h61;
	15'h2f3f: q<=8'ha5;
	15'h2f40: q<=8'h62;
	15'h2f41: q<=8'hf5;
	15'h2f42: q<=8'h90;
	15'h2f43: q<=8'h85;
	15'h2f44: q<=8'h62;
	15'h2f45: q<=8'ha5;
	15'h2f46: q<=8'h2b;
	15'h2f47: q<=8'h45;
	15'h2f48: q<=8'h9d;
	15'h2f49: q<=8'h30;
	15'h2f4a: q<=8'h0b;
	15'h2f4b: q<=8'hb9;
	15'h2f4c: q<=8'h88;
	15'h2f4d: q<=8'h00;
	15'h2f4e: q<=8'h85;
	15'h2f4f: q<=8'h63;
	15'h2f50: q<=8'hb9;
	15'h2f51: q<=8'h90;
	15'h2f52: q<=8'h00;
	15'h2f53: q<=8'hb8;
	15'h2f54: q<=8'h50;
	15'h2f55: q<=8'h11;
	15'h2f56: q<=8'hb9;
	15'h2f57: q<=8'h88;
	15'h2f58: q<=8'h00;
	15'h2f59: q<=8'h49;
	15'h2f5a: q<=8'hff;
	15'h2f5b: q<=8'h18;
	15'h2f5c: q<=8'h69;
	15'h2f5d: q<=8'h01;
	15'h2f5e: q<=8'h85;
	15'h2f5f: q<=8'h63;
	15'h2f60: q<=8'hb9;
	15'h2f61: q<=8'h90;
	15'h2f62: q<=8'h00;
	15'h2f63: q<=8'h49;
	15'h2f64: q<=8'hff;
	15'h2f65: q<=8'h69;
	15'h2f66: q<=8'h00;
	15'h2f67: q<=8'h85;
	15'h2f68: q<=8'h64;
	15'h2f69: q<=8'ha5;
	15'h2f6a: q<=8'h2d;
	15'h2f6b: q<=8'h45;
	15'h2f6c: q<=8'h9b;
	15'h2f6d: q<=8'h10;
	15'h2f6e: q<=8'h0e;
	15'h2f6f: q<=8'ha5;
	15'h2f70: q<=8'h63;
	15'h2f71: q<=8'h38;
	15'h2f72: q<=8'hf5;
	15'h2f73: q<=8'h78;
	15'h2f74: q<=8'h85;
	15'h2f75: q<=8'h63;
	15'h2f76: q<=8'ha5;
	15'h2f77: q<=8'h64;
	15'h2f78: q<=8'hf5;
	15'h2f79: q<=8'h80;
	15'h2f7a: q<=8'hb8;
	15'h2f7b: q<=8'h50;
	15'h2f7c: q<=8'h0b;
	15'h2f7d: q<=8'ha5;
	15'h2f7e: q<=8'h63;
	15'h2f7f: q<=8'h18;
	15'h2f80: q<=8'h75;
	15'h2f81: q<=8'h78;
	15'h2f82: q<=8'h85;
	15'h2f83: q<=8'h63;
	15'h2f84: q<=8'ha5;
	15'h2f85: q<=8'h64;
	15'h2f86: q<=8'h75;
	15'h2f87: q<=8'h80;
	15'h2f88: q<=8'h85;
	15'h2f89: q<=8'h64;
	15'h2f8a: q<=8'ha4;
	15'h2f8b: q<=8'ha9;
	15'h2f8c: q<=8'ha5;
	15'h2f8d: q<=8'h63;
	15'h2f8e: q<=8'h91;
	15'h2f8f: q<=8'h74;
	15'h2f90: q<=8'hc8;
	15'h2f91: q<=8'ha5;
	15'h2f92: q<=8'h64;
	15'h2f93: q<=8'h29;
	15'h2f94: q<=8'h1f;
	15'h2f95: q<=8'h91;
	15'h2f96: q<=8'h74;
	15'h2f97: q<=8'hc8;
	15'h2f98: q<=8'ha5;
	15'h2f99: q<=8'h61;
	15'h2f9a: q<=8'h91;
	15'h2f9b: q<=8'h74;
	15'h2f9c: q<=8'hc8;
	15'h2f9d: q<=8'ha5;
	15'h2f9e: q<=8'h62;
	15'h2f9f: q<=8'h29;
	15'h2fa0: q<=8'h1f;
	15'h2fa1: q<=8'h05;
	15'h2fa2: q<=8'h73;
	15'h2fa3: q<=8'h91;
	15'h2fa4: q<=8'h74;
	15'h2fa5: q<=8'hc8;
	15'h2fa6: q<=8'h84;
	15'h2fa7: q<=8'ha9;
	15'h2fa8: q<=8'hc6;
	15'h2fa9: q<=8'h99;
	15'h2faa: q<=8'hf0;
	15'h2fab: q<=8'h03;
	15'h2fac: q<=8'h4c;
	15'h2fad: q<=8'hdb;
	15'h2fae: q<=8'hbe;
	15'h2faf: q<=8'ha4;
	15'h2fb0: q<=8'ha9;
	15'h2fb1: q<=8'h88;
	15'h2fb2: q<=8'h4c;
	15'h2fb3: q<=8'h5f;
	15'h2fb4: q<=8'hdf;
	15'h2fb5: q<=8'h08;
	15'h2fb6: q<=8'h08;
	15'h2fb7: q<=8'h08;
	15'h2fb8: q<=8'h08;
	15'h2fb9: q<=8'h08;
	15'h2fba: q<=8'h08;
	15'h2fbb: q<=8'h08;
	15'h2fbc: q<=8'h08;
	15'h2fbd: q<=8'h08;
	15'h2fbe: q<=8'h09;
	15'h2fbf: q<=8'h06;
	15'h2fc0: q<=8'h07;
	15'h2fc1: q<=8'h07;
	15'h2fc2: q<=8'h04;
	15'h2fc3: q<=8'h02;
	15'h2fc4: q<=8'h00;
	15'h2fc5: q<=8'h10;
	15'h2fc6: q<=8'h20;
	15'h2fc7: q<=8'h30;
	15'h2fc8: q<=8'h40;
	15'h2fc9: q<=8'h50;
	15'h2fca: q<=8'h60;
	15'h2fcb: q<=8'h70;
	15'h2fcc: q<=8'h80;
	15'h2fcd: q<=8'h92;
	15'h2fce: q<=8'h9e;
	15'h2fcf: q<=8'hac;
	15'h2fd0: q<=8'hba;
	15'h2fd1: q<=8'hc2;
	15'h2fd2: q<=8'h0c;
	15'h2fd3: q<=8'h01;
	15'h2fd4: q<=8'h8c;
	15'h2fd5: q<=8'h01;
	15'h2fd6: q<=8'h4a;
	15'h2fd7: q<=8'h01;
	15'h2fd8: q<=8'h09;
	15'h2fd9: q<=8'h01;
	15'h2fda: q<=8'hcb;
	15'h2fdb: q<=8'h01;
	15'h2fdc: q<=8'h4b;
	15'h2fdd: q<=8'h01;
	15'h2fde: q<=8'h89;
	15'h2fdf: q<=8'h01;
	15'h2fe0: q<=8'hca;
	15'h2fe1: q<=8'h01;
	15'h2fe2: q<=8'h90;
	15'h2fe3: q<=8'h01;
	15'h2fe4: q<=8'h8a;
	15'h2fe5: q<=8'h01;
	15'h2fe6: q<=8'h23;
	15'h2fe7: q<=8'h01;
	15'h2fe8: q<=8'hdb;
	15'h2fe9: q<=8'h01;
	15'h2fea: q<=8'h41;
	15'h2feb: q<=8'h01;
	15'h2fec: q<=8'h10;
	15'h2fed: q<=8'h01;
	15'h2fee: q<=8'h0a;
	15'h2fef: q<=8'h01;
	15'h2ff0: q<=8'hcb;
	15'h2ff1: q<=8'h01;
	15'h2ff2: q<=8'h91;
	15'h2ff3: q<=8'h01;
	15'h2ff4: q<=8'h17;
	15'h2ff5: q<=8'h01;
	15'h2ff6: q<=8'h4b;
	15'h2ff7: q<=8'h01;
	15'h2ff8: q<=8'h8a;
	15'h2ff9: q<=8'h01;
	15'h2ffa: q<=8'hce;
	15'h2ffb: q<=8'h01;
	15'h2ffc: q<=8'h08;
	15'h2ffd: q<=8'h01;
	15'h2ffe: q<=8'h0a;
	15'h2fff: q<=8'h01;
	15'h3000: q<=8'hcb;
	15'h3001: q<=8'h01;
	15'h3002: q<=8'h92;
	15'h3003: q<=8'h01;
	15'h3004: q<=8'h16;
	15'h3005: q<=8'h01;
	15'h3006: q<=8'h4b;
	15'h3007: q<=8'h01;
	15'h3008: q<=8'h8a;
	15'h3009: q<=8'h01;
	15'h300a: q<=8'hcd;
	15'h300b: q<=8'h01;
	15'h300c: q<=8'h49;
	15'h300d: q<=8'h01;
	15'h300e: q<=8'h0a;
	15'h300f: q<=8'h01;
	15'h3010: q<=8'hcb;
	15'h3011: q<=8'h01;
	15'h3012: q<=8'h93;
	15'h3013: q<=8'h01;
	15'h3014: q<=8'h15;
	15'h3015: q<=8'h01;
	15'h3016: q<=8'h4b;
	15'h3017: q<=8'h01;
	15'h3018: q<=8'h8a;
	15'h3019: q<=8'h01;
	15'h301a: q<=8'hcc;
	15'h301b: q<=8'h01;
	15'h301c: q<=8'h4a;
	15'h301d: q<=8'h01;
	15'h301e: q<=8'h0a;
	15'h301f: q<=8'h01;
	15'h3020: q<=8'hcb;
	15'h3021: q<=8'h01;
	15'h3022: q<=8'h95;
	15'h3023: q<=8'h01;
	15'h3024: q<=8'h13;
	15'h3025: q<=8'h01;
	15'h3026: q<=8'h4b;
	15'h3027: q<=8'h01;
	15'h3028: q<=8'h8a;
	15'h3029: q<=8'h01;
	15'h302a: q<=8'hca;
	15'h302b: q<=8'h01;
	15'h302c: q<=8'h4c;
	15'h302d: q<=8'h01;
	15'h302e: q<=8'h0a;
	15'h302f: q<=8'h01;
	15'h3030: q<=8'hcb;
	15'h3031: q<=8'h01;
	15'h3032: q<=8'h96;
	15'h3033: q<=8'h01;
	15'h3034: q<=8'h12;
	15'h3035: q<=8'h01;
	15'h3036: q<=8'h4b;
	15'h3037: q<=8'h01;
	15'h3038: q<=8'h8a;
	15'h3039: q<=8'h01;
	15'h303a: q<=8'hc9;
	15'h303b: q<=8'h01;
	15'h303c: q<=8'h4d;
	15'h303d: q<=8'h01;
	15'h303e: q<=8'h0a;
	15'h303f: q<=8'h01;
	15'h3040: q<=8'hcb;
	15'h3041: q<=8'h01;
	15'h3042: q<=8'h97;
	15'h3043: q<=8'h01;
	15'h3044: q<=8'h11;
	15'h3045: q<=8'h01;
	15'h3046: q<=8'h4b;
	15'h3047: q<=8'h01;
	15'h3048: q<=8'h8a;
	15'h3049: q<=8'h01;
	15'h304a: q<=8'h88;
	15'h304b: q<=8'h01;
	15'h304c: q<=8'h4e;
	15'h304d: q<=8'h01;
	15'h304e: q<=8'h0a;
	15'h304f: q<=8'h01;
	15'h3050: q<=8'hcb;
	15'h3051: q<=8'h01;
	15'h3052: q<=8'h0b;
	15'h3053: q<=8'h00;
	15'h3054: q<=8'ha3;
	15'h3055: q<=8'h01;
	15'h3056: q<=8'h0a;
	15'h3057: q<=8'h01;
	15'h3058: q<=8'h10;
	15'h3059: q<=8'h01;
	15'h305a: q<=8'h4b;
	15'h305b: q<=8'h01;
	15'h305c: q<=8'h8a;
	15'h305d: q<=8'h01;
	15'h305e: q<=8'h90;
	15'h305f: q<=8'h01;
	15'h3060: q<=8'h41;
	15'h3061: q<=8'h01;
	15'h3062: q<=8'h5b;
	15'h3063: q<=8'h01;
	15'h3064: q<=8'h9a;
	15'h3065: q<=8'h01;
	15'h3066: q<=8'h31;
	15'h3067: q<=8'h01;
	15'h3068: q<=8'hb1;
	15'h3069: q<=8'h01;
	15'h306a: q<=8'h31;
	15'h306b: q<=8'h01;
	15'h306c: q<=8'hb1;
	15'h306d: q<=8'h01;
	15'h306e: q<=8'h1a;
	15'h306f: q<=8'h01;
	15'h3070: q<=8'h01;
	15'h3071: q<=8'h00;
	15'h3072: q<=8'h91;
	15'h3073: q<=8'h01;
	15'h3074: q<=8'h21;
	15'h3075: q<=8'h01;
	15'h3076: q<=8'ha1;
	15'h3077: q<=8'h01;
	15'h3078: q<=8'h21;
	15'h3079: q<=8'h01;
	15'h307a: q<=8'ha1;
	15'h307b: q<=8'h01;
	15'h307c: q<=8'h11;
	15'h307d: q<=8'h01;
	15'h307e: q<=8'h01;
	15'h307f: q<=8'h00;
	15'h3080: q<=8'h89;
	15'h3081: q<=8'h01;
	15'h3082: q<=8'h11;
	15'h3083: q<=8'h01;
	15'h3084: q<=8'h91;
	15'h3085: q<=8'h01;
	15'h3086: q<=8'h11;
	15'h3087: q<=8'h01;
	15'h3088: q<=8'h91;
	15'h3089: q<=8'h01;
	15'h308a: q<=8'h09;
	15'h308b: q<=8'h01;
	15'h308c: q<=8'h01;
	15'h308d: q<=8'h00;
	15'h308e: q<=8'h8a;
	15'h308f: q<=8'h01;
	15'h3090: q<=8'h12;
	15'h3091: q<=8'h01;
	15'h3092: q<=8'h8a;
	15'h3093: q<=8'h01;
	15'h3094: q<=8'h01;
	15'h3095: q<=8'h00;
	15'h3096: q<=8'h06;
	15'h3097: q<=8'h01;
	15'h3098: q<=8'ha5;
	15'h3099: q<=8'h57;
	15'h309a: q<=8'h38;
	15'h309b: q<=8'he5;
	15'h309c: q<=8'h5f;
	15'h309d: q<=8'h8d;
	15'h309e: q<=8'h95;
	15'h309f: q<=8'h60;
	15'h30a0: q<=8'ha9;
	15'h30a1: q<=8'h00;
	15'h30a2: q<=8'he5;
	15'h30a3: q<=8'h5b;
	15'h30a4: q<=8'h8d;
	15'h30a5: q<=8'h96;
	15'h30a6: q<=8'h60;
	15'h30a7: q<=8'h10;
	15'h30a8: q<=8'h0a;
	15'h30a9: q<=8'ha9;
	15'h30aa: q<=8'h00;
	15'h30ab: q<=8'h8d;
	15'h30ac: q<=8'h96;
	15'h30ad: q<=8'h60;
	15'h30ae: q<=8'ha9;
	15'h30af: q<=8'h01;
	15'h30b0: q<=8'h8d;
	15'h30b1: q<=8'h95;
	15'h30b2: q<=8'h60;
	15'h30b3: q<=8'ha5;
	15'h30b4: q<=8'h58;
	15'h30b5: q<=8'hc5;
	15'h30b6: q<=8'h60;
	15'h30b7: q<=8'h90;
	15'h30b8: q<=8'h07;
	15'h30b9: q<=8'he5;
	15'h30ba: q<=8'h60;
	15'h30bb: q<=8'ha2;
	15'h30bc: q<=8'h00;
	15'h30bd: q<=8'hb8;
	15'h30be: q<=8'h50;
	15'h30bf: q<=8'h07;
	15'h30c0: q<=8'ha5;
	15'h30c1: q<=8'h60;
	15'h30c2: q<=8'h38;
	15'h30c3: q<=8'he5;
	15'h30c4: q<=8'h58;
	15'h30c5: q<=8'ha2;
	15'h30c6: q<=8'hff;
	15'h30c7: q<=8'h8d;
	15'h30c8: q<=8'h8e;
	15'h30c9: q<=8'h60;
	15'h30ca: q<=8'h8d;
	15'h30cb: q<=8'h94;
	15'h30cc: q<=8'h60;
	15'h30cd: q<=8'h86;
	15'h30ce: q<=8'h33;
	15'h30cf: q<=8'ha5;
	15'h30d0: q<=8'h56;
	15'h30d1: q<=8'hc5;
	15'h30d2: q<=8'h5e;
	15'h30d3: q<=8'h90;
	15'h30d4: q<=8'h07;
	15'h30d5: q<=8'he5;
	15'h30d6: q<=8'h5e;
	15'h30d7: q<=8'ha2;
	15'h30d8: q<=8'h00;
	15'h30d9: q<=8'hb8;
	15'h30da: q<=8'h50;
	15'h30db: q<=8'h07;
	15'h30dc: q<=8'ha5;
	15'h30dd: q<=8'h5e;
	15'h30de: q<=8'h38;
	15'h30df: q<=8'he5;
	15'h30e0: q<=8'h56;
	15'h30e1: q<=8'ha2;
	15'h30e2: q<=8'hff;
	15'h30e3: q<=8'h85;
	15'h30e4: q<=8'h32;
	15'h30e5: q<=8'h86;
	15'h30e6: q<=8'h34;
	15'h30e7: q<=8'h2c;
	15'h30e8: q<=8'h40;
	15'h30e9: q<=8'h60;
	15'h30ea: q<=8'h30;
	15'h30eb: q<=8'hfb;
	15'h30ec: q<=8'had;
	15'h30ed: q<=8'h60;
	15'h30ee: q<=8'h60;
	15'h30ef: q<=8'h85;
	15'h30f0: q<=8'h63;
	15'h30f1: q<=8'had;
	15'h30f2: q<=8'h70;
	15'h30f3: q<=8'h60;
	15'h30f4: q<=8'h85;
	15'h30f5: q<=8'h64;
	15'h30f6: q<=8'ha5;
	15'h30f7: q<=8'h32;
	15'h30f8: q<=8'h8d;
	15'h30f9: q<=8'h8e;
	15'h30fa: q<=8'h60;
	15'h30fb: q<=8'h8d;
	15'h30fc: q<=8'h94;
	15'h30fd: q<=8'h60;
	15'h30fe: q<=8'ha5;
	15'h30ff: q<=8'h33;
	15'h3100: q<=8'h30;
	15'h3101: q<=8'h18;
	15'h3102: q<=8'ha5;
	15'h3103: q<=8'h63;
	15'h3104: q<=8'h18;
	15'h3105: q<=8'h65;
	15'h3106: q<=8'h68;
	15'h3107: q<=8'h85;
	15'h3108: q<=8'h63;
	15'h3109: q<=8'ha5;
	15'h310a: q<=8'h64;
	15'h310b: q<=8'h65;
	15'h310c: q<=8'h69;
	15'h310d: q<=8'h50;
	15'h310e: q<=8'h06;
	15'h310f: q<=8'ha9;
	15'h3110: q<=8'hff;
	15'h3111: q<=8'h85;
	15'h3112: q<=8'h63;
	15'h3113: q<=8'ha9;
	15'h3114: q<=8'h7f;
	15'h3115: q<=8'h85;
	15'h3116: q<=8'h64;
	15'h3117: q<=8'hb8;
	15'h3118: q<=8'h50;
	15'h3119: q<=8'h15;
	15'h311a: q<=8'ha5;
	15'h311b: q<=8'h68;
	15'h311c: q<=8'h38;
	15'h311d: q<=8'he5;
	15'h311e: q<=8'h63;
	15'h311f: q<=8'h85;
	15'h3120: q<=8'h63;
	15'h3121: q<=8'ha5;
	15'h3122: q<=8'h69;
	15'h3123: q<=8'he5;
	15'h3124: q<=8'h64;
	15'h3125: q<=8'h50;
	15'h3126: q<=8'h06;
	15'h3127: q<=8'ha9;
	15'h3128: q<=8'h00;
	15'h3129: q<=8'h85;
	15'h312a: q<=8'h63;
	15'h312b: q<=8'ha9;
	15'h312c: q<=8'h80;
	15'h312d: q<=8'h85;
	15'h312e: q<=8'h64;
	15'h312f: q<=8'h2c;
	15'h3130: q<=8'h40;
	15'h3131: q<=8'h60;
	15'h3132: q<=8'h30;
	15'h3133: q<=8'hfb;
	15'h3134: q<=8'had;
	15'h3135: q<=8'h60;
	15'h3136: q<=8'h60;
	15'h3137: q<=8'h85;
	15'h3138: q<=8'h61;
	15'h3139: q<=8'had;
	15'h313a: q<=8'h70;
	15'h313b: q<=8'h60;
	15'h313c: q<=8'h85;
	15'h313d: q<=8'h62;
	15'h313e: q<=8'ha6;
	15'h313f: q<=8'h34;
	15'h3140: q<=8'h30;
	15'h3141: q<=8'h16;
	15'h3142: q<=8'ha5;
	15'h3143: q<=8'h61;
	15'h3144: q<=8'h18;
	15'h3145: q<=8'h65;
	15'h3146: q<=8'h66;
	15'h3147: q<=8'h85;
	15'h3148: q<=8'h61;
	15'h3149: q<=8'ha5;
	15'h314a: q<=8'h62;
	15'h314b: q<=8'h65;
	15'h314c: q<=8'h67;
	15'h314d: q<=8'h50;
	15'h314e: q<=8'h06;
	15'h314f: q<=8'ha9;
	15'h3150: q<=8'hff;
	15'h3151: q<=8'h85;
	15'h3152: q<=8'h61;
	15'h3153: q<=8'ha9;
	15'h3154: q<=8'h7f;
	15'h3155: q<=8'h85;
	15'h3156: q<=8'h62;
	15'h3157: q<=8'h60;
	15'h3158: q<=8'ha5;
	15'h3159: q<=8'h66;
	15'h315a: q<=8'h38;
	15'h315b: q<=8'he5;
	15'h315c: q<=8'h61;
	15'h315d: q<=8'h85;
	15'h315e: q<=8'h61;
	15'h315f: q<=8'ha5;
	15'h3160: q<=8'h67;
	15'h3161: q<=8'he5;
	15'h3162: q<=8'h62;
	15'h3163: q<=8'h50;
	15'h3164: q<=8'h06;
	15'h3165: q<=8'ha9;
	15'h3166: q<=8'h00;
	15'h3167: q<=8'h85;
	15'h3168: q<=8'h61;
	15'h3169: q<=8'ha9;
	15'h316a: q<=8'h80;
	15'h316b: q<=8'h85;
	15'h316c: q<=8'h62;
	15'h316d: q<=8'h60;
	15'h316e: q<=8'h20;
	15'h316f: q<=8'h13;
	15'h3170: q<=8'haa;
	15'h3171: q<=8'ha9;
	15'h3172: q<=8'h80;
	15'h3173: q<=8'h85;
	15'h3174: q<=8'h5e;
	15'h3175: q<=8'ha9;
	15'h3176: q<=8'hff;
	15'h3177: q<=8'h8d;
	15'h3178: q<=8'h14;
	15'h3179: q<=8'h01;
	15'h317a: q<=8'h20;
	15'h317b: q<=8'h35;
	15'h317c: q<=8'hc2;
	15'h317d: q<=8'had;
	15'h317e: q<=8'h33;
	15'h317f: q<=8'h01;
	15'h3180: q<=8'hd0;
	15'h3181: q<=8'h03;
	15'h3182: q<=8'h8d;
	15'h3183: q<=8'h00;
	15'h3184: q<=8'h58;
	15'h3185: q<=8'ha9;
	15'h3186: q<=8'h00;
	15'h3187: q<=8'h8d;
	15'h3188: q<=8'h33;
	15'h3189: q<=8'h01;
	15'h318a: q<=8'had;
	15'h318b: q<=8'hc6;
	15'h318c: q<=8'hce;
	15'h318d: q<=8'h8d;
	15'h318e: q<=8'h00;
	15'h318f: q<=8'h20;
	15'h3190: q<=8'had;
	15'h3191: q<=8'hc7;
	15'h3192: q<=8'hce;
	15'h3193: q<=8'h8d;
	15'h3194: q<=8'h01;
	15'h3195: q<=8'h20;
	15'h3196: q<=8'ha5;
	15'h3197: q<=8'h9f;
	15'h3198: q<=8'h29;
	15'h3199: q<=8'h70;
	15'h319a: q<=8'hc9;
	15'h319b: q<=8'h5f;
	15'h319c: q<=8'h90;
	15'h319d: q<=8'h02;
	15'h319e: q<=8'ha9;
	15'h319f: q<=8'h5f;
	15'h31a0: q<=8'h4a;
	15'h31a1: q<=8'h09;
	15'h31a2: q<=8'h07;
	15'h31a3: q<=8'haa;
	15'h31a4: q<=8'ha0;
	15'h31a5: q<=8'h07;
	15'h31a6: q<=8'hbd;
	15'h31a7: q<=8'hfd;
	15'h31a8: q<=8'hc1;
	15'h31a9: q<=8'h29;
	15'h31aa: q<=8'h0f;
	15'h31ab: q<=8'h99;
	15'h31ac: q<=8'h19;
	15'h31ad: q<=8'h00;
	15'h31ae: q<=8'h99;
	15'h31af: q<=8'h00;
	15'h31b0: q<=8'h08;
	15'h31b1: q<=8'hbd;
	15'h31b2: q<=8'hfd;
	15'h31b3: q<=8'hc1;
	15'h31b4: q<=8'h4a;
	15'h31b5: q<=8'h4a;
	15'h31b6: q<=8'h4a;
	15'h31b7: q<=8'h4a;
	15'h31b8: q<=8'h99;
	15'h31b9: q<=8'h21;
	15'h31ba: q<=8'h00;
	15'h31bb: q<=8'h99;
	15'h31bc: q<=8'h08;
	15'h31bd: q<=8'h08;
	15'h31be: q<=8'hca;
	15'h31bf: q<=8'h88;
	15'h31c0: q<=8'h10;
	15'h31c1: q<=8'he4;
	15'h31c2: q<=8'h60;
	15'h31c3: q<=8'ha9;
	15'h31c4: q<=8'h00;
	15'h31c5: q<=8'h85;
	15'h31c6: q<=8'h81;
	15'h31c7: q<=8'h85;
	15'h31c8: q<=8'h91;
	15'h31c9: q<=8'h85;
	15'h31ca: q<=8'h80;
	15'h31cb: q<=8'h85;
	15'h31cc: q<=8'h78;
	15'h31cd: q<=8'h85;
	15'h31ce: q<=8'h90;
	15'h31cf: q<=8'h85;
	15'h31d0: q<=8'h88;
	15'h31d1: q<=8'ha9;
	15'h31d2: q<=8'h00;
	15'h31d3: q<=8'h8d;
	15'h31d4: q<=8'h80;
	15'h31d5: q<=8'h60;
	15'h31d6: q<=8'h8d;
	15'h31d7: q<=8'h81;
	15'h31d8: q<=8'h60;
	15'h31d9: q<=8'h8d;
	15'h31da: q<=8'h84;
	15'h31db: q<=8'h60;
	15'h31dc: q<=8'h8d;
	15'h31dd: q<=8'h85;
	15'h31de: q<=8'h60;
	15'h31df: q<=8'h8d;
	15'h31e0: q<=8'h86;
	15'h31e1: q<=8'h60;
	15'h31e2: q<=8'h8d;
	15'h31e3: q<=8'h87;
	15'h31e4: q<=8'h60;
	15'h31e5: q<=8'h8d;
	15'h31e6: q<=8'h89;
	15'h31e7: q<=8'h60;
	15'h31e8: q<=8'h8d;
	15'h31e9: q<=8'h83;
	15'h31ea: q<=8'h60;
	15'h31eb: q<=8'h8d;
	15'h31ec: q<=8'h8d;
	15'h31ed: q<=8'h60;
	15'h31ee: q<=8'h8d;
	15'h31ef: q<=8'h8e;
	15'h31f0: q<=8'h60;
	15'h31f1: q<=8'h8d;
	15'h31f2: q<=8'h8f;
	15'h31f3: q<=8'h60;
	15'h31f4: q<=8'h8d;
	15'h31f5: q<=8'h90;
	15'h31f6: q<=8'h60;
	15'h31f7: q<=8'ha9;
	15'h31f8: q<=8'h0f;
	15'h31f9: q<=8'h8d;
	15'h31fa: q<=8'h8c;
	15'h31fb: q<=8'h60;
	15'h31fc: q<=8'h60;
	15'h31fd: q<=8'h00;
	15'h31fe: q<=8'h04;
	15'h31ff: q<=8'h08;
	15'h3200: q<=8'h0c;
	15'h3201: q<=8'hc3;
	15'h3202: q<=8'h07;
	15'h3203: q<=8'h0b;
	15'h3204: q<=8'h0b;
	15'h3205: q<=8'h00;
	15'h3206: q<=8'h07;
	15'h3207: q<=8'h0b;
	15'h3208: q<=8'h08;
	15'h3209: q<=8'h44;
	15'h320a: q<=8'h03;
	15'h320b: q<=8'h0c;
	15'h320c: q<=8'h0c;
	15'h320d: q<=8'h00;
	15'h320e: q<=8'h0b;
	15'h320f: q<=8'h03;
	15'h3210: q<=8'h07;
	15'h3211: q<=8'hc8;
	15'h3212: q<=8'h0c;
	15'h3213: q<=8'h04;
	15'h3214: q<=8'h04;
	15'h3215: q<=8'h00;
	15'h3216: q<=8'h0b;
	15'h3217: q<=8'h08;
	15'h3218: q<=8'h07;
	15'h3219: q<=8'hc4;
	15'h321a: q<=8'h0c;
	15'h321b: q<=8'h03;
	15'h321c: q<=8'h03;
	15'h321d: q<=8'h00;
	15'h321e: q<=8'h04;
	15'h321f: q<=8'h08;
	15'h3220: q<=8'h0c;
	15'h3221: q<=8'hc3;
	15'h3222: q<=8'h07;
	15'h3223: q<=8'h0f;
	15'h3224: q<=8'h0b;
	15'h3225: q<=8'h00;
	15'h3226: q<=8'h0c;
	15'h3227: q<=8'h08;
	15'h3228: q<=8'h04;
	15'h3229: q<=8'hc3;
	15'h322a: q<=8'h0b;
	15'h322b: q<=8'h07;
	15'h322c: q<=8'h07;
	15'h322d: q<=8'h06;
	15'h322e: q<=8'h03;
	15'h322f: q<=8'h01;
	15'h3230: q<=8'h04;
	15'h3231: q<=8'h00;
	15'h3232: q<=8'h05;
	15'h3233: q<=8'h05;
	15'h3234: q<=8'h05;
	15'h3235: q<=8'ha6;
	15'h3236: q<=8'h3d;
	15'h3237: q<=8'hb5;
	15'h3238: q<=8'h46;
	15'h3239: q<=8'h20;
	15'h323a: q<=8'he8;
	15'h323b: q<=8'hc2;
	15'h323c: q<=8'h48;
	15'h323d: q<=8'hac;
	15'h323e: q<=8'h12;
	15'h323f: q<=8'h01;
	15'h3240: q<=8'hb9;
	15'h3241: q<=8'h8c;
	15'h3242: q<=8'hbc;
	15'h3243: q<=8'h49;
	15'h3244: q<=8'hff;
	15'h3245: q<=8'h18;
	15'h3246: q<=8'h69;
	15'h3247: q<=8'h01;
	15'h3248: q<=8'h85;
	15'h3249: q<=8'h5f;
	15'h324a: q<=8'h85;
	15'h324b: q<=8'h5d;
	15'h324c: q<=8'ha9;
	15'h324d: q<=8'h10;
	15'h324e: q<=8'h38;
	15'h324f: q<=8'he5;
	15'h3250: q<=8'h5f;
	15'h3251: q<=8'h85;
	15'h3252: q<=8'ha0;
	15'h3253: q<=8'ha9;
	15'h3254: q<=8'hff;
	15'h3255: q<=8'h85;
	15'h3256: q<=8'h5b;
	15'h3257: q<=8'hb9;
	15'h3258: q<=8'h9c;
	15'h3259: q<=8'hbc;
	15'h325a: q<=8'h85;
	15'h325b: q<=8'h60;
	15'h325c: q<=8'hb9;
	15'h325d: q<=8'hcc;
	15'h325e: q<=8'hbc;
	15'h325f: q<=8'h8d;
	15'h3260: q<=8'h11;
	15'h3261: q<=8'h01;
	15'h3262: q<=8'ha5;
	15'h3263: q<=8'h02;
	15'h3264: q<=8'hc9;
	15'h3265: q<=8'h1e;
	15'h3266: q<=8'hd0;
	15'h3267: q<=8'h0d;
	15'h3268: q<=8'hb9;
	15'h3269: q<=8'hac;
	15'h326a: q<=8'hbc;
	15'h326b: q<=8'h85;
	15'h326c: q<=8'h68;
	15'h326d: q<=8'hb9;
	15'h326e: q<=8'hbc;
	15'h326f: q<=8'hbc;
	15'h3270: q<=8'h85;
	15'h3271: q<=8'h69;
	15'h3272: q<=8'hb8;
	15'h3273: q<=8'h50;
	15'h3274: q<=8'h18;
	15'h3275: q<=8'hb9;
	15'h3276: q<=8'hac;
	15'h3277: q<=8'hbc;
	15'h3278: q<=8'h38;
	15'h3279: q<=8'he5;
	15'h327a: q<=8'h68;
	15'h327b: q<=8'h8d;
	15'h327c: q<=8'h21;
	15'h327d: q<=8'h01;
	15'h327e: q<=8'hb9;
	15'h327f: q<=8'hbc;
	15'h3280: q<=8'hbc;
	15'h3281: q<=8'hed;
	15'h3282: q<=8'h69;
	15'h3283: q<=8'h00;
	15'h3284: q<=8'ha2;
	15'h3285: q<=8'h03;
	15'h3286: q<=8'h4a;
	15'h3287: q<=8'h6e;
	15'h3288: q<=8'h21;
	15'h3289: q<=8'h01;
	15'h328a: q<=8'hca;
	15'h328b: q<=8'h10;
	15'h328c: q<=8'hf9;
	15'h328d: q<=8'ha9;
	15'h328e: q<=8'h00;
	15'h328f: q<=8'h85;
	15'h3290: q<=8'h66;
	15'h3291: q<=8'h85;
	15'h3292: q<=8'h67;
	15'h3293: q<=8'ha9;
	15'h3294: q<=8'h00;
	15'h3295: q<=8'h8d;
	15'h3296: q<=8'h0f;
	15'h3297: q<=8'h01;
	15'h3298: q<=8'h8d;
	15'h3299: q<=8'h10;
	15'h329a: q<=8'h01;
	15'h329b: q<=8'ha9;
	15'h329c: q<=8'h2c;
	15'h329d: q<=8'h8d;
	15'h329e: q<=8'h13;
	15'h329f: q<=8'h01;
	15'h32a0: q<=8'h68;
	15'h32a1: q<=8'ha8;
	15'h32a2: q<=8'ha2;
	15'h32a3: q<=8'h0f;
	15'h32a4: q<=8'hb9;
	15'h32a5: q<=8'h7c;
	15'h32a6: q<=8'hb9;
	15'h32a7: q<=8'h9d;
	15'h32a8: q<=8'hce;
	15'h32a9: q<=8'h03;
	15'h32aa: q<=8'hb9;
	15'h32ab: q<=8'h7c;
	15'h32ac: q<=8'hba;
	15'h32ad: q<=8'h9d;
	15'h32ae: q<=8'hde;
	15'h32af: q<=8'h03;
	15'h32b0: q<=8'ha9;
	15'h32b1: q<=8'h00;
	15'h32b2: q<=8'h9d;
	15'h32b3: q<=8'h1a;
	15'h32b4: q<=8'h03;
	15'h32b5: q<=8'h9d;
	15'h32b6: q<=8'h3a;
	15'h32b7: q<=8'h03;
	15'h32b8: q<=8'h9d;
	15'h32b9: q<=8'h9a;
	15'h32ba: q<=8'h03;
	15'h32bb: q<=8'hb9;
	15'h32bc: q<=8'h7c;
	15'h32bd: q<=8'hbb;
	15'h32be: q<=8'h9d;
	15'h32bf: q<=8'hee;
	15'h32c0: q<=8'h03;
	15'h32c1: q<=8'h88;
	15'h32c2: q<=8'hca;
	15'h32c3: q<=8'h10;
	15'h32c4: q<=8'hdf;
	15'h32c5: q<=8'ha0;
	15'h32c6: q<=8'h00;
	15'h32c7: q<=8'ha2;
	15'h32c8: q<=8'h0f;
	15'h32c9: q<=8'hb9;
	15'h32ca: q<=8'hce;
	15'h32cb: q<=8'h03;
	15'h32cc: q<=8'h38;
	15'h32cd: q<=8'h7d;
	15'h32ce: q<=8'hce;
	15'h32cf: q<=8'h03;
	15'h32d0: q<=8'h6a;
	15'h32d1: q<=8'h9d;
	15'h32d2: q<=8'h35;
	15'h32d3: q<=8'h04;
	15'h32d4: q<=8'hb9;
	15'h32d5: q<=8'hde;
	15'h32d6: q<=8'h03;
	15'h32d7: q<=8'h38;
	15'h32d8: q<=8'h7d;
	15'h32d9: q<=8'hde;
	15'h32da: q<=8'h03;
	15'h32db: q<=8'h6a;
	15'h32dc: q<=8'h9d;
	15'h32dd: q<=8'h45;
	15'h32de: q<=8'h04;
	15'h32df: q<=8'h88;
	15'h32e0: q<=8'h10;
	15'h32e1: q<=8'h02;
	15'h32e2: q<=8'ha0;
	15'h32e3: q<=8'h0f;
	15'h32e4: q<=8'hca;
	15'h32e5: q<=8'h10;
	15'h32e6: q<=8'he2;
	15'h32e7: q<=8'h60;
	15'h32e8: q<=8'ha2;
	15'h32e9: q<=8'h00;
	15'h32ea: q<=8'hc9;
	15'h32eb: q<=8'h62;
	15'h32ec: q<=8'h90;
	15'h32ed: q<=8'h05;
	15'h32ee: q<=8'had;
	15'h32ef: q<=8'hca;
	15'h32f0: q<=8'h60;
	15'h32f1: q<=8'h29;
	15'h32f2: q<=8'h5f;
	15'h32f3: q<=8'hc9;
	15'h32f4: q<=8'h10;
	15'h32f5: q<=8'h90;
	15'h32f6: q<=8'h04;
	15'h32f7: q<=8'he8;
	15'h32f8: q<=8'h38;
	15'h32f9: q<=8'he9;
	15'h32fa: q<=8'h10;
	15'h32fb: q<=8'hc9;
	15'h32fc: q<=8'h10;
	15'h32fd: q<=8'hb0;
	15'h32fe: q<=8'hf6;
	15'h32ff: q<=8'ha8;
	15'h3300: q<=8'hb9;
	15'h3301: q<=8'h7c;
	15'h3302: q<=8'hbc;
	15'h3303: q<=8'h8d;
	15'h3304: q<=8'h12;
	15'h3305: q<=8'h01;
	15'h3306: q<=8'h0a;
	15'h3307: q<=8'h0a;
	15'h3308: q<=8'h0a;
	15'h3309: q<=8'h0a;
	15'h330a: q<=8'h09;
	15'h330b: q<=8'h0f;
	15'h330c: q<=8'h60;
	15'h330d: q<=8'had;
	15'h330e: q<=8'h10;
	15'h330f: q<=8'h01;
	15'h3310: q<=8'hd0;
	15'h3311: q<=8'h27;
	15'h3312: q<=8'ha9;
	15'h3313: q<=8'hf0;
	15'h3314: q<=8'h85;
	15'h3315: q<=8'h57;
	15'h3316: q<=8'ha2;
	15'h3317: q<=8'h4f;
	15'h3318: q<=8'h20;
	15'h3319: q<=8'h73;
	15'h331a: q<=8'hc4;
	15'h331b: q<=8'h8d;
	15'h331c: q<=8'h10;
	15'h331d: q<=8'h01;
	15'h331e: q<=8'hf0;
	15'h331f: q<=8'h03;
	15'h3320: q<=8'h8d;
	15'h3321: q<=8'h0f;
	15'h3322: q<=8'h01;
	15'h3323: q<=8'had;
	15'h3324: q<=8'h0f;
	15'h3325: q<=8'h01;
	15'h3326: q<=8'hd0;
	15'h3327: q<=8'h11;
	15'h3328: q<=8'ha9;
	15'h3329: q<=8'h10;
	15'h332a: q<=8'h85;
	15'h332b: q<=8'h57;
	15'h332c: q<=8'h20;
	15'h332d: q<=8'h53;
	15'h332e: q<=8'hc4;
	15'h332f: q<=8'ha5;
	15'h3330: q<=8'h57;
	15'h3331: q<=8'ha2;
	15'h3332: q<=8'h0f;
	15'h3333: q<=8'h20;
	15'h3334: q<=8'h73;
	15'h3335: q<=8'hc4;
	15'h3336: q<=8'h8d;
	15'h3337: q<=8'h0f;
	15'h3338: q<=8'h01;
	15'h3339: q<=8'ha9;
	15'h333a: q<=8'h01;
	15'h333b: q<=8'h20;
	15'h333c: q<=8'h6a;
	15'h333d: q<=8'hdf;
	15'h333e: q<=8'ha0;
	15'h333f: q<=8'h06;
	15'h3340: q<=8'h84;
	15'h3341: q<=8'h9e;
	15'h3342: q<=8'hae;
	15'h3343: q<=8'h10;
	15'h3344: q<=8'h01;
	15'h3345: q<=8'hf0;
	15'h3346: q<=8'h01;
	15'h3347: q<=8'h60;
	15'h3348: q<=8'hae;
	15'h3349: q<=8'h13;
	15'h334a: q<=8'h01;
	15'h334b: q<=8'hd0;
	15'h334c: q<=8'h01;
	15'h334d: q<=8'h60;
	15'h334e: q<=8'ha2;
	15'h334f: q<=8'h0f;
	15'h3350: q<=8'ha9;
	15'h3351: q<=8'hc0;
	15'h3352: q<=8'h20;
	15'h3353: q<=8'hee;
	15'h3354: q<=8'hc3;
	15'h3355: q<=8'hca;
	15'h3356: q<=8'h10;
	15'h3357: q<=8'hf8;
	15'h3358: q<=8'ha0;
	15'h3359: q<=8'h06;
	15'h335a: q<=8'h84;
	15'h335b: q<=8'h9e;
	15'h335c: q<=8'ha9;
	15'h335d: q<=8'h08;
	15'h335e: q<=8'h20;
	15'h335f: q<=8'h4c;
	15'h3360: q<=8'hdf;
	15'h3361: q<=8'ha0;
	15'h3362: q<=8'h4f;
	15'h3363: q<=8'had;
	15'h3364: q<=8'h10;
	15'h3365: q<=8'h01;
	15'h3366: q<=8'h20;
	15'h3367: q<=8'h6e;
	15'h3368: q<=8'hc3;
	15'h3369: q<=8'ha0;
	15'h336a: q<=8'h0f;
	15'h336b: q<=8'had;
	15'h336c: q<=8'h0f;
	15'h336d: q<=8'h01;
	15'h336e: q<=8'hd0;
	15'h336f: q<=8'h49;
	15'h3370: q<=8'h84;
	15'h3371: q<=8'h37;
	15'h3372: q<=8'hb9;
	15'h3373: q<=8'h2a;
	15'h3374: q<=8'h03;
	15'h3375: q<=8'h85;
	15'h3376: q<=8'h61;
	15'h3377: q<=8'hb9;
	15'h3378: q<=8'h1a;
	15'h3379: q<=8'h03;
	15'h337a: q<=8'h85;
	15'h337b: q<=8'h62;
	15'h337c: q<=8'hb9;
	15'h337d: q<=8'h4a;
	15'h337e: q<=8'h03;
	15'h337f: q<=8'h85;
	15'h3380: q<=8'h63;
	15'h3381: q<=8'hb9;
	15'h3382: q<=8'h3a;
	15'h3383: q<=8'h03;
	15'h3384: q<=8'h85;
	15'h3385: q<=8'h64;
	15'h3386: q<=8'ha2;
	15'h3387: q<=8'h61;
	15'h3388: q<=8'h20;
	15'h3389: q<=8'h72;
	15'h338a: q<=8'hc7;
	15'h338b: q<=8'ha5;
	15'h338c: q<=8'h74;
	15'h338d: q<=8'h85;
	15'h338e: q<=8'hb0;
	15'h338f: q<=8'ha5;
	15'h3390: q<=8'h75;
	15'h3391: q<=8'h85;
	15'h3392: q<=8'hb1;
	15'h3393: q<=8'ha2;
	15'h3394: q<=8'h0f;
	15'h3395: q<=8'had;
	15'h3396: q<=8'h11;
	15'h3397: q<=8'h01;
	15'h3398: q<=8'hf0;
	15'h3399: q<=8'h01;
	15'h339a: q<=8'hca;
	15'h339b: q<=8'ha9;
	15'h339c: q<=8'hc0;
	15'h339d: q<=8'h85;
	15'h339e: q<=8'h73;
	15'h339f: q<=8'h86;
	15'h33a0: q<=8'h38;
	15'h33a1: q<=8'hc6;
	15'h33a2: q<=8'h37;
	15'h33a3: q<=8'ha5;
	15'h33a4: q<=8'h37;
	15'h33a5: q<=8'h29;
	15'h33a6: q<=8'h0f;
	15'h33a7: q<=8'hc9;
	15'h33a8: q<=8'h0f;
	15'h33a9: q<=8'hd0;
	15'h33aa: q<=8'h07;
	15'h33ab: q<=8'ha5;
	15'h33ac: q<=8'h37;
	15'h33ad: q<=8'h18;
	15'h33ae: q<=8'h69;
	15'h33af: q<=8'h10;
	15'h33b0: q<=8'h85;
	15'h33b1: q<=8'h37;
	15'h33b2: q<=8'h20;
	15'h33b3: q<=8'h23;
	15'h33b4: q<=8'hc4;
	15'h33b5: q<=8'hc6;
	15'h33b6: q<=8'h38;
	15'h33b7: q<=8'h10;
	15'h33b8: q<=8'he8;
	15'h33b9: q<=8'h60;
	15'h33ba: q<=8'ha5;
	15'h33bb: q<=8'h61;
	15'h33bc: q<=8'h38;
	15'h33bd: q<=8'he5;
	15'h33be: q<=8'h6a;
	15'h33bf: q<=8'h85;
	15'h33c0: q<=8'h6e;
	15'h33c1: q<=8'ha5;
	15'h33c2: q<=8'h62;
	15'h33c3: q<=8'he5;
	15'h33c4: q<=8'h6b;
	15'h33c5: q<=8'h85;
	15'h33c6: q<=8'h6f;
	15'h33c7: q<=8'ha5;
	15'h33c8: q<=8'h63;
	15'h33c9: q<=8'h38;
	15'h33ca: q<=8'he5;
	15'h33cb: q<=8'h6c;
	15'h33cc: q<=8'h85;
	15'h33cd: q<=8'h70;
	15'h33ce: q<=8'ha5;
	15'h33cf: q<=8'h64;
	15'h33d0: q<=8'he5;
	15'h33d1: q<=8'h6d;
	15'h33d2: q<=8'h85;
	15'h33d3: q<=8'h71;
	15'h33d4: q<=8'ha2;
	15'h33d5: q<=8'h6e;
	15'h33d6: q<=8'h20;
	15'h33d7: q<=8'h92;
	15'h33d8: q<=8'hdf;
	15'h33d9: q<=8'ha5;
	15'h33da: q<=8'h61;
	15'h33db: q<=8'h85;
	15'h33dc: q<=8'h6a;
	15'h33dd: q<=8'ha5;
	15'h33de: q<=8'h62;
	15'h33df: q<=8'h85;
	15'h33e0: q<=8'h6b;
	15'h33e1: q<=8'ha5;
	15'h33e2: q<=8'h63;
	15'h33e3: q<=8'h85;
	15'h33e4: q<=8'h6c;
	15'h33e5: q<=8'ha5;
	15'h33e6: q<=8'h64;
	15'h33e7: q<=8'h85;
	15'h33e8: q<=8'h6d;
	15'h33e9: q<=8'ha9;
	15'h33ea: q<=8'hc0;
	15'h33eb: q<=8'h85;
	15'h33ec: q<=8'h73;
	15'h33ed: q<=8'h60;
	15'h33ee: q<=8'h86;
	15'h33ef: q<=8'h37;
	15'h33f0: q<=8'h48;
	15'h33f1: q<=8'ha4;
	15'h33f2: q<=8'h9e;
	15'h33f3: q<=8'ha9;
	15'h33f4: q<=8'h08;
	15'h33f5: q<=8'h20;
	15'h33f6: q<=8'h4c;
	15'h33f7: q<=8'hdf;
	15'h33f8: q<=8'h20;
	15'h33f9: q<=8'h3c;
	15'h33fa: q<=8'hc4;
	15'h33fb: q<=8'ha2;
	15'h33fc: q<=8'h61;
	15'h33fd: q<=8'h20;
	15'h33fe: q<=8'h72;
	15'h33ff: q<=8'hc7;
	15'h3400: q<=8'h68;
	15'h3401: q<=8'h85;
	15'h3402: q<=8'h73;
	15'h3403: q<=8'h48;
	15'h3404: q<=8'h20;
	15'h3405: q<=8'h23;
	15'h3406: q<=8'hc4;
	15'h3407: q<=8'hc6;
	15'h3408: q<=8'h37;
	15'h3409: q<=8'ha4;
	15'h340a: q<=8'h9e;
	15'h340b: q<=8'ha9;
	15'h340c: q<=8'h00;
	15'h340d: q<=8'h85;
	15'h340e: q<=8'h73;
	15'h340f: q<=8'ha9;
	15'h3410: q<=8'h08;
	15'h3411: q<=8'h20;
	15'h3412: q<=8'h4c;
	15'h3413: q<=8'hdf;
	15'h3414: q<=8'h20;
	15'h3415: q<=8'h23;
	15'h3416: q<=8'hc4;
	15'h3417: q<=8'h68;
	15'h3418: q<=8'h85;
	15'h3419: q<=8'h73;
	15'h341a: q<=8'h20;
	15'h341b: q<=8'h3c;
	15'h341c: q<=8'hc4;
	15'h341d: q<=8'h20;
	15'h341e: q<=8'hba;
	15'h341f: q<=8'hc3;
	15'h3420: q<=8'ha6;
	15'h3421: q<=8'h37;
	15'h3422: q<=8'h60;
	15'h3423: q<=8'ha6;
	15'h3424: q<=8'h37;
	15'h3425: q<=8'hbd;
	15'h3426: q<=8'h2a;
	15'h3427: q<=8'h03;
	15'h3428: q<=8'h85;
	15'h3429: q<=8'h61;
	15'h342a: q<=8'hbd;
	15'h342b: q<=8'h1a;
	15'h342c: q<=8'h03;
	15'h342d: q<=8'h85;
	15'h342e: q<=8'h62;
	15'h342f: q<=8'hbd;
	15'h3430: q<=8'h4a;
	15'h3431: q<=8'h03;
	15'h3432: q<=8'h85;
	15'h3433: q<=8'h63;
	15'h3434: q<=8'hbd;
	15'h3435: q<=8'h3a;
	15'h3436: q<=8'h03;
	15'h3437: q<=8'h85;
	15'h3438: q<=8'h64;
	15'h3439: q<=8'h4c;
	15'h343a: q<=8'hba;
	15'h343b: q<=8'hc3;
	15'h343c: q<=8'ha6;
	15'h343d: q<=8'h37;
	15'h343e: q<=8'hbd;
	15'h343f: q<=8'h6a;
	15'h3440: q<=8'h03;
	15'h3441: q<=8'h85;
	15'h3442: q<=8'h61;
	15'h3443: q<=8'hbd;
	15'h3444: q<=8'h5a;
	15'h3445: q<=8'h03;
	15'h3446: q<=8'h85;
	15'h3447: q<=8'h62;
	15'h3448: q<=8'hbd;
	15'h3449: q<=8'h8a;
	15'h344a: q<=8'h03;
	15'h344b: q<=8'h85;
	15'h344c: q<=8'h63;
	15'h344d: q<=8'hbd;
	15'h344e: q<=8'h7a;
	15'h344f: q<=8'h03;
	15'h3450: q<=8'h85;
	15'h3451: q<=8'h64;
	15'h3452: q<=8'h60;
	15'h3453: q<=8'ha5;
	15'h3454: q<=8'h5b;
	15'h3455: q<=8'hd0;
	15'h3456: q<=8'h1a;
	15'h3457: q<=8'ha5;
	15'h3458: q<=8'h57;
	15'h3459: q<=8'h38;
	15'h345a: q<=8'he5;
	15'h345b: q<=8'h5f;
	15'h345c: q<=8'h90;
	15'h345d: q<=8'h02;
	15'h345e: q<=8'hc9;
	15'h345f: q<=8'h0c;
	15'h3460: q<=8'hb0;
	15'h3461: q<=8'h0f;
	15'h3462: q<=8'ha5;
	15'h3463: q<=8'h5f;
	15'h3464: q<=8'h18;
	15'h3465: q<=8'h69;
	15'h3466: q<=8'h0f;
	15'h3467: q<=8'hb0;
	15'h3468: q<=8'h02;
	15'h3469: q<=8'hc9;
	15'h346a: q<=8'hf0;
	15'h346b: q<=8'h90;
	15'h346c: q<=8'h02;
	15'h346d: q<=8'ha9;
	15'h346e: q<=8'hf0;
	15'h346f: q<=8'h85;
	15'h3470: q<=8'h57;
	15'h3471: q<=8'h60;
	15'h3472: q<=8'hdb;
	15'h3473: q<=8'h85;
	15'h3474: q<=8'h57;
	15'h3475: q<=8'h86;
	15'h3476: q<=8'h38;
	15'h3477: q<=8'ha9;
	15'h3478: q<=8'h00;
	15'h3479: q<=8'h85;
	15'h347a: q<=8'h59;
	15'h347b: q<=8'ha2;
	15'h347c: q<=8'h0f;
	15'h347d: q<=8'h86;
	15'h347e: q<=8'h37;
	15'h347f: q<=8'ha6;
	15'h3480: q<=8'h37;
	15'h3481: q<=8'hbd;
	15'h3482: q<=8'hce;
	15'h3483: q<=8'h03;
	15'h3484: q<=8'h85;
	15'h3485: q<=8'h56;
	15'h3486: q<=8'hbd;
	15'h3487: q<=8'hde;
	15'h3488: q<=8'h03;
	15'h3489: q<=8'h85;
	15'h348a: q<=8'h58;
	15'h348b: q<=8'h20;
	15'h348c: q<=8'h98;
	15'h348d: q<=8'hc0;
	15'h348e: q<=8'ha6;
	15'h348f: q<=8'h38;
	15'h3490: q<=8'ha4;
	15'h3491: q<=8'h61;
	15'h3492: q<=8'ha5;
	15'h3493: q<=8'h62;
	15'h3494: q<=8'h30;
	15'h3495: q<=8'h0d;
	15'h3496: q<=8'hc9;
	15'h3497: q<=8'h04;
	15'h3498: q<=8'h90;
	15'h3499: q<=8'h06;
	15'h349a: q<=8'ha0;
	15'h349b: q<=8'hff;
	15'h349c: q<=8'ha9;
	15'h349d: q<=8'h03;
	15'h349e: q<=8'he6;
	15'h349f: q<=8'h59;
	15'h34a0: q<=8'hb8;
	15'h34a1: q<=8'h50;
	15'h34a2: q<=8'h0a;
	15'h34a3: q<=8'hc9;
	15'h34a4: q<=8'hfc;
	15'h34a5: q<=8'hb0;
	15'h34a6: q<=8'h06;
	15'h34a7: q<=8'ha0;
	15'h34a8: q<=8'h01;
	15'h34a9: q<=8'ha9;
	15'h34aa: q<=8'hfc;
	15'h34ab: q<=8'he6;
	15'h34ac: q<=8'h59;
	15'h34ad: q<=8'h9d;
	15'h34ae: q<=8'h1a;
	15'h34af: q<=8'h03;
	15'h34b0: q<=8'h98;
	15'h34b1: q<=8'h9d;
	15'h34b2: q<=8'h2a;
	15'h34b3: q<=8'h03;
	15'h34b4: q<=8'ha4;
	15'h34b5: q<=8'h63;
	15'h34b6: q<=8'ha5;
	15'h34b7: q<=8'h64;
	15'h34b8: q<=8'h30;
	15'h34b9: q<=8'h0d;
	15'h34ba: q<=8'hc9;
	15'h34bb: q<=8'h04;
	15'h34bc: q<=8'h90;
	15'h34bd: q<=8'h06;
	15'h34be: q<=8'ha0;
	15'h34bf: q<=8'hff;
	15'h34c0: q<=8'ha9;
	15'h34c1: q<=8'h03;
	15'h34c2: q<=8'he6;
	15'h34c3: q<=8'h59;
	15'h34c4: q<=8'hb8;
	15'h34c5: q<=8'h50;
	15'h34c6: q<=8'h0a;
	15'h34c7: q<=8'hc9;
	15'h34c8: q<=8'hfc;
	15'h34c9: q<=8'hb0;
	15'h34ca: q<=8'h06;
	15'h34cb: q<=8'ha9;
	15'h34cc: q<=8'hfc;
	15'h34cd: q<=8'ha0;
	15'h34ce: q<=8'h01;
	15'h34cf: q<=8'he6;
	15'h34d0: q<=8'h59;
	15'h34d1: q<=8'h9d;
	15'h34d2: q<=8'h3a;
	15'h34d3: q<=8'h03;
	15'h34d4: q<=8'h98;
	15'h34d5: q<=8'h9d;
	15'h34d6: q<=8'h4a;
	15'h34d7: q<=8'h03;
	15'h34d8: q<=8'hc6;
	15'h34d9: q<=8'h38;
	15'h34da: q<=8'hc6;
	15'h34db: q<=8'h37;
	15'h34dc: q<=8'h10;
	15'h34dd: q<=8'ha1;
	15'h34de: q<=8'ha5;
	15'h34df: q<=8'h59;
	15'h34e0: q<=8'h60;
	15'h34e1: q<=8'h20;
	15'h34e2: q<=8'he8;
	15'h34e3: q<=8'hc2;
	15'h34e4: q<=8'h85;
	15'h34e5: q<=8'h36;
	15'h34e6: q<=8'h86;
	15'h34e7: q<=8'h35;
	15'h34e8: q<=8'ha9;
	15'h34e9: q<=8'h00;
	15'h34ea: q<=8'h85;
	15'h34eb: q<=8'h73;
	15'h34ec: q<=8'ha9;
	15'h34ed: q<=8'h05;
	15'h34ee: q<=8'h20;
	15'h34ef: q<=8'h6a;
	15'h34f0: q<=8'hdf;
	15'h34f1: q<=8'ha5;
	15'h34f2: q<=8'h35;
	15'h34f3: q<=8'h29;
	15'h34f4: q<=8'h07;
	15'h34f5: q<=8'haa;
	15'h34f6: q<=8'hbc;
	15'h34f7: q<=8'h2d;
	15'h34f8: q<=8'hc2;
	15'h34f9: q<=8'h84;
	15'h34fa: q<=8'h9e;
	15'h34fb: q<=8'ha9;
	15'h34fc: q<=8'h08;
	15'h34fd: q<=8'h20;
	15'h34fe: q<=8'h4c;
	15'h34ff: q<=8'hdf;
	15'h3500: q<=8'hae;
	15'h3501: q<=8'h12;
	15'h3502: q<=8'h01;
	15'h3503: q<=8'ha5;
	15'h3504: q<=8'h36;
	15'h3505: q<=8'hbc;
	15'h3506: q<=8'hcc;
	15'h3507: q<=8'hbc;
	15'h3508: q<=8'hd0;
	15'h3509: q<=8'h03;
	15'h350a: q<=8'h38;
	15'h350b: q<=8'he9;
	15'h350c: q<=8'h0f;
	15'h350d: q<=8'ha8;
	15'h350e: q<=8'hb9;
	15'h350f: q<=8'h7c;
	15'h3510: q<=8'hba;
	15'h3511: q<=8'h85;
	15'h3512: q<=8'h57;
	15'h3513: q<=8'h49;
	15'h3514: q<=8'h80;
	15'h3515: q<=8'haa;
	15'h3516: q<=8'hb9;
	15'h3517: q<=8'h7c;
	15'h3518: q<=8'hb9;
	15'h3519: q<=8'h85;
	15'h351a: q<=8'h56;
	15'h351b: q<=8'h49;
	15'h351c: q<=8'h80;
	15'h351d: q<=8'h20;
	15'h351e: q<=8'h75;
	15'h351f: q<=8'hdf;
	15'h3520: q<=8'ha9;
	15'h3521: q<=8'hc0;
	15'h3522: q<=8'h85;
	15'h3523: q<=8'h73;
	15'h3524: q<=8'ha2;
	15'h3525: q<=8'h0f;
	15'h3526: q<=8'h86;
	15'h3527: q<=8'h38;
	15'h3528: q<=8'ha4;
	15'h3529: q<=8'h36;
	15'h352a: q<=8'hb9;
	15'h352b: q<=8'h7c;
	15'h352c: q<=8'hb9;
	15'h352d: q<=8'haa;
	15'h352e: q<=8'h38;
	15'h352f: q<=8'he5;
	15'h3530: q<=8'h56;
	15'h3531: q<=8'h48;
	15'h3532: q<=8'h86;
	15'h3533: q<=8'h56;
	15'h3534: q<=8'hb9;
	15'h3535: q<=8'h7c;
	15'h3536: q<=8'hba;
	15'h3537: q<=8'ha8;
	15'h3538: q<=8'h38;
	15'h3539: q<=8'he5;
	15'h353a: q<=8'h57;
	15'h353b: q<=8'haa;
	15'h353c: q<=8'h84;
	15'h353d: q<=8'h57;
	15'h353e: q<=8'h68;
	15'h353f: q<=8'h20;
	15'h3540: q<=8'h75;
	15'h3541: q<=8'hdf;
	15'h3542: q<=8'hc6;
	15'h3543: q<=8'h36;
	15'h3544: q<=8'hc6;
	15'h3545: q<=8'h38;
	15'h3546: q<=8'h10;
	15'h3547: q<=8'he0;
	15'h3548: q<=8'ha9;
	15'h3549: q<=8'h01;
	15'h354a: q<=8'h4c;
	15'h354b: q<=8'h6a;
	15'h354c: q<=8'hdf;
	15'h354d: q<=8'had;
	15'h354e: q<=8'h15;
	15'h354f: q<=8'h01;
	15'h3550: q<=8'hf0;
	15'h3551: q<=8'h5f;
	15'h3552: q<=8'ha5;
	15'h3553: q<=8'h5f;
	15'h3554: q<=8'h48;
	15'h3555: q<=8'ha5;
	15'h3556: q<=8'h5b;
	15'h3557: q<=8'h48;
	15'h3558: q<=8'ha5;
	15'h3559: q<=8'ha0;
	15'h355a: q<=8'h48;
	15'h355b: q<=8'ha9;
	15'h355c: q<=8'he8;
	15'h355d: q<=8'h85;
	15'h355e: q<=8'h5f;
	15'h355f: q<=8'ha9;
	15'h3560: q<=8'hff;
	15'h3561: q<=8'h85;
	15'h3562: q<=8'h5b;
	15'h3563: q<=8'ha9;
	15'h3564: q<=8'h28;
	15'h3565: q<=8'h85;
	15'h3566: q<=8'ha0;
	15'h3567: q<=8'ha2;
	15'h3568: q<=8'h07;
	15'h3569: q<=8'h86;
	15'h356a: q<=8'h37;
	15'h356b: q<=8'ha6;
	15'h356c: q<=8'h37;
	15'h356d: q<=8'hbd;
	15'h356e: q<=8'hfe;
	15'h356f: q<=8'h03;
	15'h3570: q<=8'hf0;
	15'h3571: q<=8'h32;
	15'h3572: q<=8'h85;
	15'h3573: q<=8'h57;
	15'h3574: q<=8'ha9;
	15'h3575: q<=8'h80;
	15'h3576: q<=8'h85;
	15'h3577: q<=8'h56;
	15'h3578: q<=8'ha9;
	15'h3579: q<=8'h80;
	15'h357a: q<=8'h85;
	15'h357b: q<=8'h58;
	15'h357c: q<=8'ha5;
	15'h357d: q<=8'h9f;
	15'h357e: q<=8'hc9;
	15'h357f: q<=8'h05;
	15'h3580: q<=8'hb0;
	15'h3581: q<=8'h05;
	15'h3582: q<=8'ha9;
	15'h3583: q<=8'h06;
	15'h3584: q<=8'hb8;
	15'h3585: q<=8'h50;
	15'h3586: q<=8'h09;
	15'h3587: q<=8'h8a;
	15'h3588: q<=8'h29;
	15'h3589: q<=8'h07;
	15'h358a: q<=8'hc9;
	15'h358b: q<=8'h07;
	15'h358c: q<=8'hd0;
	15'h358d: q<=8'h02;
	15'h358e: q<=8'ha9;
	15'h358f: q<=8'h04;
	15'h3590: q<=8'h85;
	15'h3591: q<=8'h9e;
	15'h3592: q<=8'ha8;
	15'h3593: q<=8'ha9;
	15'h3594: q<=8'h08;
	15'h3595: q<=8'h20;
	15'h3596: q<=8'h4c;
	15'h3597: q<=8'hdf;
	15'h3598: q<=8'ha5;
	15'h3599: q<=8'h37;
	15'h359a: q<=8'h29;
	15'h359b: q<=8'h03;
	15'h359c: q<=8'h0a;
	15'h359d: q<=8'h69;
	15'h359e: q<=8'h0a;
	15'h359f: q<=8'h85;
	15'h35a0: q<=8'h55;
	15'h35a1: q<=8'h20;
	15'h35a2: q<=8'h09;
	15'h35a3: q<=8'hbd;
	15'h35a4: q<=8'hc6;
	15'h35a5: q<=8'h37;
	15'h35a6: q<=8'h10;
	15'h35a7: q<=8'hc3;
	15'h35a8: q<=8'h68;
	15'h35a9: q<=8'h85;
	15'h35aa: q<=8'ha0;
	15'h35ab: q<=8'h68;
	15'h35ac: q<=8'h85;
	15'h35ad: q<=8'h5b;
	15'h35ae: q<=8'h68;
	15'h35af: q<=8'h85;
	15'h35b0: q<=8'h5f;
	15'h35b1: q<=8'had;
	15'h35b2: q<=8'h1f;
	15'h35b3: q<=8'h01;
	15'h35b4: q<=8'hf0;
	15'h35b5: q<=8'h0b;
	15'h35b6: q<=8'ha6;
	15'h35b7: q<=8'h42;
	15'h35b8: q<=8'he0;
	15'h35b9: q<=8'h15;
	15'h35ba: q<=8'h90;
	15'h35bb: q<=8'h05;
	15'h35bc: q<=8'ha6;
	15'h35bd: q<=8'h40;
	15'h35be: q<=8'hfe;
	15'h35bf: q<=8'h00;
	15'h35c0: q<=8'h02;
	15'h35c1: q<=8'h60;
	15'h35c2: q<=8'had;
	15'h35c3: q<=8'h10;
	15'h35c4: q<=8'h01;
	15'h35c5: q<=8'hf0;
	15'h35c6: q<=8'h01;
	15'h35c7: q<=8'h60;
	15'h35c8: q<=8'ha5;
	15'h35c9: q<=8'h5b;
	15'h35ca: q<=8'hd0;
	15'h35cb: q<=8'h07;
	15'h35cc: q<=8'ha5;
	15'h35cd: q<=8'h5f;
	15'h35ce: q<=8'hc9;
	15'h35cf: q<=8'hf0;
	15'h35d0: q<=8'h90;
	15'h35d1: q<=8'h01;
	15'h35d2: q<=8'h60;
	15'h35d3: q<=8'ha9;
	15'h35d4: q<=8'h01;
	15'h35d5: q<=8'h20;
	15'h35d6: q<=8'h6a;
	15'h35d7: q<=8'hdf;
	15'h35d8: q<=8'ha5;
	15'h35d9: q<=8'h74;
	15'h35da: q<=8'h48;
	15'h35db: q<=8'ha5;
	15'h35dc: q<=8'h75;
	15'h35dd: q<=8'h48;
	15'h35de: q<=8'ha9;
	15'h35df: q<=8'h00;
	15'h35e0: q<=8'h85;
	15'h35e1: q<=8'h38;
	15'h35e2: q<=8'h85;
	15'h35e3: q<=8'ha9;
	15'h35e4: q<=8'ha2;
	15'h35e5: q<=8'h0f;
	15'h35e6: q<=8'had;
	15'h35e7: q<=8'h11;
	15'h35e8: q<=8'h01;
	15'h35e9: q<=8'hf0;
	15'h35ea: q<=8'h01;
	15'h35eb: q<=8'hca;
	15'h35ec: q<=8'h86;
	15'h35ed: q<=8'h37;
	15'h35ee: q<=8'ha2;
	15'h35ef: q<=8'h03;
	15'h35f0: q<=8'ha4;
	15'h35f1: q<=8'ha9;
	15'h35f2: q<=8'hbd;
	15'h35f3: q<=8'h69;
	15'h35f4: q<=8'hc6;
	15'h35f5: q<=8'h91;
	15'h35f6: q<=8'h74;
	15'h35f7: q<=8'hc8;
	15'h35f8: q<=8'hca;
	15'h35f9: q<=8'h10;
	15'h35fa: q<=8'hf7;
	15'h35fb: q<=8'h84;
	15'h35fc: q<=8'ha9;
	15'h35fd: q<=8'had;
	15'h35fe: q<=8'h14;
	15'h35ff: q<=8'h01;
	15'h3600: q<=8'hd0;
	15'h3601: q<=8'h4a;
	15'h3602: q<=8'ha6;
	15'h3603: q<=8'h38;
	15'h3604: q<=8'hbd;
	15'h3605: q<=8'h9a;
	15'h3606: q<=8'h03;
	15'h3607: q<=8'h30;
	15'h3608: q<=8'h11;
	15'h3609: q<=8'ha2;
	15'h360a: q<=8'h0b;
	15'h360b: q<=8'ha4;
	15'h360c: q<=8'ha9;
	15'h360d: q<=8'hb1;
	15'h360e: q<=8'haa;
	15'h360f: q<=8'h91;
	15'h3610: q<=8'h74;
	15'h3611: q<=8'hc8;
	15'h3612: q<=8'hca;
	15'h3613: q<=8'h10;
	15'h3614: q<=8'hf8;
	15'h3615: q<=8'h84;
	15'h3616: q<=8'ha9;
	15'h3617: q<=8'hb8;
	15'h3618: q<=8'h50;
	15'h3619: q<=8'h2f;
	15'h361a: q<=8'ha4;
	15'h361b: q<=8'ha9;
	15'h361c: q<=8'hb1;
	15'h361d: q<=8'haa;
	15'h361e: q<=8'h91;
	15'h361f: q<=8'h74;
	15'h3620: q<=8'h85;
	15'h3621: q<=8'h6c;
	15'h3622: q<=8'hc8;
	15'h3623: q<=8'hb1;
	15'h3624: q<=8'haa;
	15'h3625: q<=8'h91;
	15'h3626: q<=8'h74;
	15'h3627: q<=8'hc9;
	15'h3628: q<=8'h10;
	15'h3629: q<=8'h90;
	15'h362a: q<=8'h02;
	15'h362b: q<=8'h09;
	15'h362c: q<=8'he0;
	15'h362d: q<=8'h85;
	15'h362e: q<=8'h6d;
	15'h362f: q<=8'hc8;
	15'h3630: q<=8'hb1;
	15'h3631: q<=8'haa;
	15'h3632: q<=8'h91;
	15'h3633: q<=8'h74;
	15'h3634: q<=8'h85;
	15'h3635: q<=8'h6a;
	15'h3636: q<=8'hc8;
	15'h3637: q<=8'hb1;
	15'h3638: q<=8'haa;
	15'h3639: q<=8'h91;
	15'h363a: q<=8'h74;
	15'h363b: q<=8'hc9;
	15'h363c: q<=8'h10;
	15'h363d: q<=8'h90;
	15'h363e: q<=8'h02;
	15'h363f: q<=8'h09;
	15'h3640: q<=8'he0;
	15'h3641: q<=8'h85;
	15'h3642: q<=8'h6b;
	15'h3643: q<=8'hc8;
	15'h3644: q<=8'h84;
	15'h3645: q<=8'ha9;
	15'h3646: q<=8'h20;
	15'h3647: q<=8'hc7;
	15'h3648: q<=8'hc6;
	15'h3649: q<=8'hb8;
	15'h364a: q<=8'h50;
	15'h364b: q<=8'h06;
	15'h364c: q<=8'h20;
	15'h364d: q<=8'h6d;
	15'h364e: q<=8'hc6;
	15'h364f: q<=8'h20;
	15'h3650: q<=8'hc7;
	15'h3651: q<=8'hc6;
	15'h3652: q<=8'ha6;
	15'h3653: q<=8'h38;
	15'h3654: q<=8'h1e;
	15'h3655: q<=8'h9a;
	15'h3656: q<=8'h03;
	15'h3657: q<=8'he6;
	15'h3658: q<=8'h38;
	15'h3659: q<=8'hc6;
	15'h365a: q<=8'h37;
	15'h365b: q<=8'h10;
	15'h365c: q<=8'h91;
	15'h365d: q<=8'h68;
	15'h365e: q<=8'h85;
	15'h365f: q<=8'hab;
	15'h3660: q<=8'h68;
	15'h3661: q<=8'h85;
	15'h3662: q<=8'haa;
	15'h3663: q<=8'ha4;
	15'h3664: q<=8'ha9;
	15'h3665: q<=8'h88;
	15'h3666: q<=8'h4c;
	15'h3667: q<=8'h5f;
	15'h3668: q<=8'hdf;
	15'h3669: q<=8'h80;
	15'h366a: q<=8'h40;
	15'h366b: q<=8'h68;
	15'h366c: q<=8'h05;
	15'h366d: q<=8'ha5;
	15'h366e: q<=8'h38;
	15'h366f: q<=8'haa;
	15'h3670: q<=8'h18;
	15'h3671: q<=8'h69;
	15'h3672: q<=8'h01;
	15'h3673: q<=8'h29;
	15'h3674: q<=8'h0f;
	15'h3675: q<=8'ha8;
	15'h3676: q<=8'hbd;
	15'h3677: q<=8'h6a;
	15'h3678: q<=8'h03;
	15'h3679: q<=8'h38;
	15'h367a: q<=8'h79;
	15'h367b: q<=8'h6a;
	15'h367c: q<=8'h03;
	15'h367d: q<=8'h85;
	15'h367e: q<=8'h61;
	15'h367f: q<=8'hbd;
	15'h3680: q<=8'h5a;
	15'h3681: q<=8'h03;
	15'h3682: q<=8'h79;
	15'h3683: q<=8'h5a;
	15'h3684: q<=8'h03;
	15'h3685: q<=8'h85;
	15'h3686: q<=8'h62;
	15'h3687: q<=8'h0a;
	15'h3688: q<=8'h66;
	15'h3689: q<=8'h62;
	15'h368a: q<=8'h66;
	15'h368b: q<=8'h61;
	15'h368c: q<=8'hbd;
	15'h368d: q<=8'h8a;
	15'h368e: q<=8'h03;
	15'h368f: q<=8'h38;
	15'h3690: q<=8'h79;
	15'h3691: q<=8'h8a;
	15'h3692: q<=8'h03;
	15'h3693: q<=8'h85;
	15'h3694: q<=8'h63;
	15'h3695: q<=8'hbd;
	15'h3696: q<=8'h7a;
	15'h3697: q<=8'h03;
	15'h3698: q<=8'h79;
	15'h3699: q<=8'h7a;
	15'h369a: q<=8'h03;
	15'h369b: q<=8'h85;
	15'h369c: q<=8'h64;
	15'h369d: q<=8'h0a;
	15'h369e: q<=8'h66;
	15'h369f: q<=8'h64;
	15'h36a0: q<=8'h66;
	15'h36a1: q<=8'h63;
	15'h36a2: q<=8'ha4;
	15'h36a3: q<=8'ha9;
	15'h36a4: q<=8'ha5;
	15'h36a5: q<=8'h63;
	15'h36a6: q<=8'h91;
	15'h36a7: q<=8'h74;
	15'h36a8: q<=8'hc8;
	15'h36a9: q<=8'h85;
	15'h36aa: q<=8'h6c;
	15'h36ab: q<=8'ha5;
	15'h36ac: q<=8'h64;
	15'h36ad: q<=8'h85;
	15'h36ae: q<=8'h6d;
	15'h36af: q<=8'h29;
	15'h36b0: q<=8'h1f;
	15'h36b1: q<=8'h91;
	15'h36b2: q<=8'h74;
	15'h36b3: q<=8'hc8;
	15'h36b4: q<=8'ha5;
	15'h36b5: q<=8'h61;
	15'h36b6: q<=8'h91;
	15'h36b7: q<=8'h74;
	15'h36b8: q<=8'hc8;
	15'h36b9: q<=8'h85;
	15'h36ba: q<=8'h6a;
	15'h36bb: q<=8'ha5;
	15'h36bc: q<=8'h62;
	15'h36bd: q<=8'h85;
	15'h36be: q<=8'h6b;
	15'h36bf: q<=8'h29;
	15'h36c0: q<=8'h1f;
	15'h36c1: q<=8'h91;
	15'h36c2: q<=8'h74;
	15'h36c3: q<=8'hc8;
	15'h36c4: q<=8'h84;
	15'h36c5: q<=8'ha9;
	15'h36c6: q<=8'h60;
	15'h36c7: q<=8'ha6;
	15'h36c8: q<=8'h38;
	15'h36c9: q<=8'hbd;
	15'h36ca: q<=8'hac;
	15'h36cb: q<=8'h03;
	15'h36cc: q<=8'hd0;
	15'h36cd: q<=8'h16;
	15'h36ce: q<=8'ha4;
	15'h36cf: q<=8'ha9;
	15'h36d0: q<=8'ha2;
	15'h36d1: q<=8'h03;
	15'h36d2: q<=8'ha9;
	15'h36d3: q<=8'h00;
	15'h36d4: q<=8'h91;
	15'h36d5: q<=8'h74;
	15'h36d6: q<=8'hc8;
	15'h36d7: q<=8'ha9;
	15'h36d8: q<=8'h71;
	15'h36d9: q<=8'h91;
	15'h36da: q<=8'h74;
	15'h36db: q<=8'hc8;
	15'h36dc: q<=8'hca;
	15'h36dd: q<=8'h10;
	15'h36de: q<=8'hf3;
	15'h36df: q<=8'h84;
	15'h36e0: q<=8'ha9;
	15'h36e1: q<=8'hb8;
	15'h36e2: q<=8'h50;
	15'h36e3: q<=8'h57;
	15'h36e4: q<=8'h85;
	15'h36e5: q<=8'h57;
	15'h36e6: q<=8'h20;
	15'h36e7: q<=8'h53;
	15'h36e8: q<=8'hc4;
	15'h36e9: q<=8'hbd;
	15'h36ea: q<=8'h35;
	15'h36eb: q<=8'h04;
	15'h36ec: q<=8'h85;
	15'h36ed: q<=8'h56;
	15'h36ee: q<=8'hbd;
	15'h36ef: q<=8'h45;
	15'h36f0: q<=8'h04;
	15'h36f1: q<=8'h85;
	15'h36f2: q<=8'h58;
	15'h36f3: q<=8'h20;
	15'h36f4: q<=8'h98;
	15'h36f5: q<=8'hc0;
	15'h36f6: q<=8'h20;
	15'h36f7: q<=8'h3c;
	15'h36f8: q<=8'hc7;
	15'h36f9: q<=8'ha6;
	15'h36fa: q<=8'h38;
	15'h36fb: q<=8'hbd;
	15'h36fc: q<=8'h9a;
	15'h36fd: q<=8'h03;
	15'h36fe: q<=8'h29;
	15'h36ff: q<=8'h40;
	15'h3700: q<=8'hf0;
	15'h3701: q<=8'h1f;
	15'h3702: q<=8'h20;
	15'h3703: q<=8'h3e;
	15'h3704: q<=8'hbd;
	15'h3705: q<=8'had;
	15'h3706: q<=8'hca;
	15'h3707: q<=8'h60;
	15'h3708: q<=8'h29;
	15'h3709: q<=8'h02;
	15'h370a: q<=8'h18;
	15'h370b: q<=8'h69;
	15'h370c: q<=8'h1c;
	15'h370d: q<=8'haa;
	15'h370e: q<=8'hbd;
	15'h370f: q<=8'hc9;
	15'h3710: q<=8'hce;
	15'h3711: q<=8'hc8;
	15'h3712: q<=8'h91;
	15'h3713: q<=8'h74;
	15'h3714: q<=8'h88;
	15'h3715: q<=8'hbd;
	15'h3716: q<=8'hc8;
	15'h3717: q<=8'hce;
	15'h3718: q<=8'h91;
	15'h3719: q<=8'h74;
	15'h371a: q<=8'hc8;
	15'h371b: q<=8'hc8;
	15'h371c: q<=8'h84;
	15'h371d: q<=8'ha9;
	15'h371e: q<=8'hb8;
	15'h371f: q<=8'h50;
	15'h3720: q<=8'h1a;
	15'h3721: q<=8'ha4;
	15'h3722: q<=8'ha9;
	15'h3723: q<=8'ha9;
	15'h3724: q<=8'h00;
	15'h3725: q<=8'h91;
	15'h3726: q<=8'h74;
	15'h3727: q<=8'hc8;
	15'h3728: q<=8'ha9;
	15'h3729: q<=8'h68;
	15'h372a: q<=8'h91;
	15'h372b: q<=8'h74;
	15'h372c: q<=8'hc8;
	15'h372d: q<=8'had;
	15'h372e: q<=8'hb2;
	15'h372f: q<=8'h3d;
	15'h3730: q<=8'h91;
	15'h3731: q<=8'h74;
	15'h3732: q<=8'hc8;
	15'h3733: q<=8'had;
	15'h3734: q<=8'hb3;
	15'h3735: q<=8'h3d;
	15'h3736: q<=8'h91;
	15'h3737: q<=8'h74;
	15'h3738: q<=8'hc8;
	15'h3739: q<=8'h84;
	15'h373a: q<=8'ha9;
	15'h373b: q<=8'h60;
	15'h373c: q<=8'ha4;
	15'h373d: q<=8'ha9;
	15'h373e: q<=8'ha5;
	15'h373f: q<=8'h63;
	15'h3740: q<=8'h38;
	15'h3741: q<=8'he5;
	15'h3742: q<=8'h6c;
	15'h3743: q<=8'h91;
	15'h3744: q<=8'h74;
	15'h3745: q<=8'hc8;
	15'h3746: q<=8'ha5;
	15'h3747: q<=8'h64;
	15'h3748: q<=8'he5;
	15'h3749: q<=8'h6d;
	15'h374a: q<=8'h29;
	15'h374b: q<=8'h1f;
	15'h374c: q<=8'h91;
	15'h374d: q<=8'h74;
	15'h374e: q<=8'hc8;
	15'h374f: q<=8'ha5;
	15'h3750: q<=8'h61;
	15'h3751: q<=8'h38;
	15'h3752: q<=8'he5;
	15'h3753: q<=8'h6a;
	15'h3754: q<=8'h91;
	15'h3755: q<=8'h74;
	15'h3756: q<=8'hc8;
	15'h3757: q<=8'ha5;
	15'h3758: q<=8'h62;
	15'h3759: q<=8'he5;
	15'h375a: q<=8'h6b;
	15'h375b: q<=8'h29;
	15'h375c: q<=8'h1f;
	15'h375d: q<=8'h09;
	15'h375e: q<=8'ha0;
	15'h375f: q<=8'h91;
	15'h3760: q<=8'h74;
	15'h3761: q<=8'hc8;
	15'h3762: q<=8'h84;
	15'h3763: q<=8'ha9;
	15'h3764: q<=8'h60;
	15'h3765: q<=8'ha0;
	15'h3766: q<=8'h00;
	15'h3767: q<=8'h98;
	15'h3768: q<=8'h91;
	15'h3769: q<=8'h74;
	15'h376a: q<=8'ha9;
	15'h376b: q<=8'h71;
	15'h376c: q<=8'hc8;
	15'h376d: q<=8'h91;
	15'h376e: q<=8'h74;
	15'h376f: q<=8'hc8;
	15'h3770: q<=8'hd0;
	15'h3771: q<=8'h02;
	15'h3772: q<=8'ha0;
	15'h3773: q<=8'h00;
	15'h3774: q<=8'ha9;
	15'h3775: q<=8'h40;
	15'h3776: q<=8'h91;
	15'h3777: q<=8'h74;
	15'h3778: q<=8'ha9;
	15'h3779: q<=8'h80;
	15'h377a: q<=8'hc8;
	15'h377b: q<=8'h91;
	15'h377c: q<=8'h74;
	15'h377d: q<=8'hc8;
	15'h377e: q<=8'hb5;
	15'h377f: q<=8'h02;
	15'h3780: q<=8'h85;
	15'h3781: q<=8'h6c;
	15'h3782: q<=8'h91;
	15'h3783: q<=8'h74;
	15'h3784: q<=8'hc8;
	15'h3785: q<=8'hb5;
	15'h3786: q<=8'h03;
	15'h3787: q<=8'h85;
	15'h3788: q<=8'h6d;
	15'h3789: q<=8'h29;
	15'h378a: q<=8'h1f;
	15'h378b: q<=8'h91;
	15'h378c: q<=8'h74;
	15'h378d: q<=8'hb5;
	15'h378e: q<=8'h00;
	15'h378f: q<=8'h85;
	15'h3790: q<=8'h6a;
	15'h3791: q<=8'hc8;
	15'h3792: q<=8'h91;
	15'h3793: q<=8'h74;
	15'h3794: q<=8'hb5;
	15'h3795: q<=8'h01;
	15'h3796: q<=8'h85;
	15'h3797: q<=8'h6b;
	15'h3798: q<=8'h29;
	15'h3799: q<=8'h1f;
	15'h379a: q<=8'hc8;
	15'h379b: q<=8'h91;
	15'h379c: q<=8'h74;
	15'h379d: q<=8'h4c;
	15'h379e: q<=8'h5f;
	15'h379f: q<=8'hdf;
	15'h37a0: q<=8'h20;
	15'h37a1: q<=8'h95;
	15'h37a2: q<=8'hcd;
	15'h37a3: q<=8'ha9;
	15'h37a4: q<=8'h00;
	15'h37a5: q<=8'h85;
	15'h37a6: q<=8'h00;
	15'h37a7: q<=8'ha5;
	15'h37a8: q<=8'h53;
	15'h37a9: q<=8'hc9;
	15'h37aa: q<=8'h09;
	15'h37ab: q<=8'h90;
	15'h37ac: q<=8'hfa;
	15'h37ad: q<=8'ha9;
	15'h37ae: q<=8'h00;
	15'h37af: q<=8'h85;
	15'h37b0: q<=8'h53;
	15'h37b1: q<=8'h20;
	15'h37b2: q<=8'hbd;
	15'h37b3: q<=8'hc7;
	15'h37b4: q<=8'h20;
	15'h37b5: q<=8'h91;
	15'h37b6: q<=8'hc8;
	15'h37b7: q<=8'h20;
	15'h37b8: q<=8'hb6;
	15'h37b9: q<=8'hb1;
	15'h37ba: q<=8'h18;
	15'h37bb: q<=8'h90;
	15'h37bc: q<=8'hea;
	15'h37bd: q<=8'had;
	15'h37be: q<=8'h00;
	15'h37bf: q<=8'h0d;
	15'h37c0: q<=8'h29;
	15'h37c1: q<=8'h83;
	15'h37c2: q<=8'hc9;
	15'h37c3: q<=8'h82;
	15'h37c4: q<=8'hf0;
	15'h37c5: q<=8'h13;
	15'h37c6: q<=8'h20;
	15'h37c7: q<=8'hd2;
	15'h37c8: q<=8'ha7;
	15'h37c9: q<=8'ha6;
	15'h37ca: q<=8'h00;
	15'h37cb: q<=8'ha5;
	15'h37cc: q<=8'h4e;
	15'h37cd: q<=8'h09;
	15'h37ce: q<=8'h80;
	15'h37cf: q<=8'h85;
	15'h37d0: q<=8'h4e;
	15'h37d1: q<=8'hbd;
	15'h37d2: q<=8'hdb;
	15'h37d3: q<=8'hc7;
	15'h37d4: q<=8'h48;
	15'h37d5: q<=8'hbd;
	15'h37d6: q<=8'hda;
	15'h37d7: q<=8'hc7;
	15'h37d8: q<=8'h48;
	15'h37d9: q<=8'h60;
	15'h37da: q<=8'h0b;
	15'h37db: q<=8'hc9;
	15'h37dc: q<=8'h3f;
	15'h37dd: q<=8'hc9;
	15'h37de: q<=8'h0a;
	15'h37df: q<=8'h97;
	15'h37e0: q<=8'hae;
	15'h37e1: q<=8'hc9;
	15'h37e2: q<=8'hf0;
	15'h37e3: q<=8'hc9;
	15'h37e4: q<=8'hff;
	15'h37e5: q<=8'hc7;
	15'h37e6: q<=8'h00;
	15'h37e7: q<=8'h00;
	15'h37e8: q<=8'h8b;
	15'h37e9: q<=8'hc9;
	15'h37ea: q<=8'h3e;
	15'h37eb: q<=8'hac;
	15'h37ec: q<=8'h6d;
	15'h37ed: q<=8'had;
	15'h37ee: q<=8'h17;
	15'h37ef: q<=8'hca;
	15'h37f0: q<=8'h48;
	15'h37f1: q<=8'h91;
	15'h37f2: q<=8'h4a;
	15'h37f3: q<=8'h90;
	15'h37f4: q<=8'he6;
	15'h37f5: q<=8'hb0;
	15'h37f6: q<=8'h07;
	15'h37f7: q<=8'h91;
	15'h37f8: q<=8'h7a;
	15'h37f9: q<=8'hc9;
	15'h37fa: q<=8'h28;
	15'h37fb: q<=8'h97;
	15'h37fc: q<=8'he0;
	15'h37fd: q<=8'hd7;
	15'h37fe: q<=8'h17;
	15'h37ff: q<=8'ha6;
	15'h3800: q<=8'ha5;
	15'h3801: q<=8'h03;
	15'h3802: q<=8'h2d;
	15'h3803: q<=8'h6b;
	15'h3804: q<=8'h01;
	15'h3805: q<=8'hd0;
	15'h3806: q<=8'h11;
	15'h3807: q<=8'ha5;
	15'h3808: q<=8'h04;
	15'h3809: q<=8'hf0;
	15'h380a: q<=8'h02;
	15'h380b: q<=8'hc6;
	15'h380c: q<=8'h04;
	15'h380d: q<=8'hd0;
	15'h380e: q<=8'h09;
	15'h380f: q<=8'ha5;
	15'h3810: q<=8'h02;
	15'h3811: q<=8'h85;
	15'h3812: q<=8'h00;
	15'h3813: q<=8'ha9;
	15'h3814: q<=8'h00;
	15'h3815: q<=8'h8d;
	15'h3816: q<=8'h6b;
	15'h3817: q<=8'h01;
	15'h3818: q<=8'h4c;
	15'h3819: q<=8'h49;
	15'h381a: q<=8'h97;
	15'h381b: q<=8'ha5;
	15'h381c: q<=8'h06;
	15'h381d: q<=8'ha0;
	15'h381e: q<=8'h00;
	15'h381f: q<=8'hc9;
	15'h3820: q<=8'h02;
	15'h3821: q<=8'ha5;
	15'h3822: q<=8'h4e;
	15'h3823: q<=8'h29;
	15'h3824: q<=8'h60;
	15'h3825: q<=8'h84;
	15'h3826: q<=8'h4e;
	15'h3827: q<=8'hf0;
	15'h3828: q<=8'h48;
	15'h3829: q<=8'hb0;
	15'h382a: q<=8'h05;
	15'h382b: q<=8'h29;
	15'h382c: q<=8'h20;
	15'h382d: q<=8'hb8;
	15'h382e: q<=8'h50;
	15'h382f: q<=8'h05;
	15'h3830: q<=8'hc8;
	15'h3831: q<=8'hc6;
	15'h3832: q<=8'h06;
	15'h3833: q<=8'h29;
	15'h3834: q<=8'h40;
	15'h3835: q<=8'hf0;
	15'h3836: q<=8'h03;
	15'h3837: q<=8'hc6;
	15'h3838: q<=8'h06;
	15'h3839: q<=8'hc8;
	15'h383a: q<=8'h98;
	15'h383b: q<=8'h85;
	15'h383c: q<=8'h3e;
	15'h383d: q<=8'hf0;
	15'h383e: q<=8'h2f;
	15'h383f: q<=8'ha5;
	15'h3840: q<=8'h05;
	15'h3841: q<=8'h09;
	15'h3842: q<=8'hc0;
	15'h3843: q<=8'h85;
	15'h3844: q<=8'h05;
	15'h3845: q<=8'ha9;
	15'h3846: q<=8'h00;
	15'h3847: q<=8'h85;
	15'h3848: q<=8'h16;
	15'h3849: q<=8'h85;
	15'h384a: q<=8'h18;
	15'h384b: q<=8'ha9;
	15'h384c: q<=8'h00;
	15'h384d: q<=8'h85;
	15'h384e: q<=8'h00;
	15'h384f: q<=8'hc6;
	15'h3850: q<=8'h3e;
	15'h3851: q<=8'ha6;
	15'h3852: q<=8'h3e;
	15'h3853: q<=8'hf0;
	15'h3854: q<=8'h02;
	15'h3855: q<=8'ha2;
	15'h3856: q<=8'h03;
	15'h3857: q<=8'hfe;
	15'h3858: q<=8'h0c;
	15'h3859: q<=8'h04;
	15'h385a: q<=8'hd0;
	15'h385b: q<=8'h03;
	15'h385c: q<=8'hfe;
	15'h385d: q<=8'h0d;
	15'h385e: q<=8'h04;
	15'h385f: q<=8'had;
	15'h3860: q<=8'h00;
	15'h3861: q<=8'h01;
	15'h3862: q<=8'h38;
	15'h3863: q<=8'h65;
	15'h3864: q<=8'h3e;
	15'h3865: q<=8'hc9;
	15'h3866: q<=8'h63;
	15'h3867: q<=8'h90;
	15'h3868: q<=8'h02;
	15'h3869: q<=8'ha9;
	15'h386a: q<=8'h63;
	15'h386b: q<=8'h8d;
	15'h386c: q<=8'h00;
	15'h386d: q<=8'h01;
	15'h386e: q<=8'hb8;
	15'h386f: q<=8'h50;
	15'h3870: q<=8'h1f;
	15'h3871: q<=8'ha5;
	15'h3872: q<=8'h50;
	15'h3873: q<=8'hf0;
	15'h3874: q<=8'h1b;
	15'h3875: q<=8'h24;
	15'h3876: q<=8'h05;
	15'h3877: q<=8'h30;
	15'h3878: q<=8'h17;
	15'h3879: q<=8'ha9;
	15'h387a: q<=8'h10;
	15'h387b: q<=8'h85;
	15'h387c: q<=8'h01;
	15'h387d: q<=8'ha9;
	15'h387e: q<=8'h20;
	15'h387f: q<=8'h85;
	15'h3880: q<=8'h04;
	15'h3881: q<=8'ha9;
	15'h3882: q<=8'h0a;
	15'h3883: q<=8'h85;
	15'h3884: q<=8'h00;
	15'h3885: q<=8'ha9;
	15'h3886: q<=8'h14;
	15'h3887: q<=8'h85;
	15'h3888: q<=8'h02;
	15'h3889: q<=8'ha9;
	15'h388a: q<=8'h00;
	15'h388b: q<=8'h85;
	15'h388c: q<=8'h50;
	15'h388d: q<=8'h8d;
	15'h388e: q<=8'h23;
	15'h388f: q<=8'h01;
	15'h3890: q<=8'h60;
	15'h3891: q<=8'had;
	15'h3892: q<=8'h00;
	15'h3893: q<=8'h0c;
	15'h3894: q<=8'h29;
	15'h3895: q<=8'h10;
	15'h3896: q<=8'hd0;
	15'h3897: q<=8'h07;
	15'h3898: q<=8'ha9;
	15'h3899: q<=8'h22;
	15'h389a: q<=8'h85;
	15'h389b: q<=8'h00;
	15'h389c: q<=8'hb8;
	15'h389d: q<=8'h50;
	15'h389e: q<=8'h44;
	15'h389f: q<=8'h24;
	15'h38a0: q<=8'h05;
	15'h38a1: q<=8'h70;
	15'h38a2: q<=8'h40;
	15'h38a3: q<=8'ha5;
	15'h38a4: q<=8'h0a;
	15'h38a5: q<=8'h29;
	15'h38a6: q<=8'h01;
	15'h38a7: q<=8'hf0;
	15'h38a8: q<=8'h29;
	15'h38a9: q<=8'ha4;
	15'h38aa: q<=8'h06;
	15'h38ab: q<=8'hd0;
	15'h38ac: q<=8'h04;
	15'h38ad: q<=8'ha9;
	15'h38ae: q<=8'h80;
	15'h38af: q<=8'h85;
	15'h38b0: q<=8'ha2;
	15'h38b1: q<=8'h24;
	15'h38b2: q<=8'ha2;
	15'h38b3: q<=8'h10;
	15'h38b4: q<=8'h1d;
	15'h38b5: q<=8'hc0;
	15'h38b6: q<=8'h02;
	15'h38b7: q<=8'hb0;
	15'h38b8: q<=8'h11;
	15'h38b9: q<=8'h98;
	15'h38ba: q<=8'hf0;
	15'h38bb: q<=8'h08;
	15'h38bc: q<=8'ha9;
	15'h38bd: q<=8'h16;
	15'h38be: q<=8'h85;
	15'h38bf: q<=8'h01;
	15'h38c0: q<=8'ha9;
	15'h38c1: q<=8'h0a;
	15'h38c2: q<=8'h85;
	15'h38c3: q<=8'h00;
	15'h38c4: q<=8'h4c;
	15'h38c5: q<=8'hd9;
	15'h38c6: q<=8'hc8;
	15'h38c7: q<=8'hb8;
	15'h38c8: q<=8'h50;
	15'h38c9: q<=8'h08;
	15'h38ca: q<=8'ha9;
	15'h38cb: q<=8'h14;
	15'h38cc: q<=8'h85;
	15'h38cd: q<=8'h00;
	15'h38ce: q<=8'ha9;
	15'h38cf: q<=8'h00;
	15'h38d0: q<=8'h85;
	15'h38d1: q<=8'ha2;
	15'h38d2: q<=8'ha5;
	15'h38d3: q<=8'h06;
	15'h38d4: q<=8'hf0;
	15'h38d5: q<=8'h03;
	15'h38d6: q<=8'h20;
	15'h38d7: q<=8'h1b;
	15'h38d8: q<=8'hc8;
	15'h38d9: q<=8'ha5;
	15'h38da: q<=8'h09;
	15'h38db: q<=8'h29;
	15'h38dc: q<=8'h03;
	15'h38dd: q<=8'hd0;
	15'h38de: q<=8'h04;
	15'h38df: q<=8'ha9;
	15'h38e0: q<=8'h02;
	15'h38e1: q<=8'h85;
	15'h38e2: q<=8'h06;
	15'h38e3: q<=8'he6;
	15'h38e4: q<=8'h03;
	15'h38e5: q<=8'ha5;
	15'h38e6: q<=8'h03;
	15'h38e7: q<=8'h29;
	15'h38e8: q<=8'h01;
	15'h38e9: q<=8'hf0;
	15'h38ea: q<=8'h03;
	15'h38eb: q<=8'h20;
	15'h38ec: q<=8'h1b;
	15'h38ed: q<=8'hde;
	15'h38ee: q<=8'ha5;
	15'h38ef: q<=8'h0c;
	15'h38f0: q<=8'hf0;
	15'h38f1: q<=8'h03;
	15'h38f2: q<=8'h20;
	15'h38f3: q<=8'hfa;
	15'h38f4: q<=8'hcc;
	15'h38f5: q<=8'had;
	15'h38f6: q<=8'h6c;
	15'h38f7: q<=8'h01;
	15'h38f8: q<=8'hf0;
	15'h38f9: q<=8'h07;
	15'h38fa: q<=8'ha9;
	15'h38fb: q<=8'h13;
	15'h38fc: q<=8'hc5;
	15'h38fd: q<=8'h9f;
	15'h38fe: q<=8'hb0;
	15'h38ff: q<=8'h01;
	15'h3900: q<=8'hf8;
	15'h3901: q<=8'ha5;
	15'h3902: q<=8'h4e;
	15'h3903: q<=8'h29;
	15'h3904: q<=8'h80;
	15'h3905: q<=8'hf0;
	15'h3906: q<=8'h04;
	15'h3907: q<=8'ha9;
	15'h3908: q<=8'h00;
	15'h3909: q<=8'h85;
	15'h390a: q<=8'h4e;
	15'h390b: q<=8'h60;
	15'h390c: q<=8'h20;
	15'h390d: q<=8'ha2;
	15'h390e: q<=8'hab;
	15'h390f: q<=8'h20;
	15'h3910: q<=8'h6e;
	15'h3911: q<=8'hc1;
	15'h3912: q<=8'ha5;
	15'h3913: q<=8'h05;
	15'h3914: q<=8'h10;
	15'h3915: q<=8'h03;
	15'h3916: q<=8'h20;
	15'h3917: q<=8'h62;
	15'h3918: q<=8'hca;
	15'h3919: q<=8'ha9;
	15'h391a: q<=8'h00;
	15'h391b: q<=8'h85;
	15'h391c: q<=8'h49;
	15'h391d: q<=8'ha6;
	15'h391e: q<=8'h3e;
	15'h391f: q<=8'h86;
	15'h3920: q<=8'h3d;
	15'h3921: q<=8'ha6;
	15'h3922: q<=8'h3d;
	15'h3923: q<=8'had;
	15'h3924: q<=8'h58;
	15'h3925: q<=8'h01;
	15'h3926: q<=8'h9d;
	15'h3927: q<=8'h48;
	15'h3928: q<=8'h00;
	15'h3929: q<=8'ha9;
	15'h392a: q<=8'hff;
	15'h392b: q<=8'h9d;
	15'h392c: q<=8'h46;
	15'h392d: q<=8'h00;
	15'h392e: q<=8'hc6;
	15'h392f: q<=8'h3d;
	15'h3930: q<=8'h10;
	15'h3931: q<=8'hef;
	15'h3932: q<=8'ha9;
	15'h3933: q<=8'h00;
	15'h3934: q<=8'h85;
	15'h3935: q<=8'h3f;
	15'h3936: q<=8'h8d;
	15'h3937: q<=8'h15;
	15'h3938: q<=8'h01;
	15'h3939: q<=8'ha5;
	15'h393a: q<=8'h3e;
	15'h393b: q<=8'h85;
	15'h393c: q<=8'h3d;
	15'h393d: q<=8'h4c;
	15'h393e: q<=8'hc4;
	15'h393f: q<=8'h90;
	15'h3940: q<=8'ha9;
	15'h3941: q<=8'h00;
	15'h3942: q<=8'h85;
	15'h3943: q<=8'h01;
	15'h3944: q<=8'ha9;
	15'h3945: q<=8'h1e;
	15'h3946: q<=8'h85;
	15'h3947: q<=8'h00;
	15'h3948: q<=8'h85;
	15'h3949: q<=8'h02;
	15'h394a: q<=8'ha5;
	15'h394b: q<=8'h3f;
	15'h394c: q<=8'hc5;
	15'h394d: q<=8'h3d;
	15'h394e: q<=8'hf0;
	15'h394f: q<=8'h1c;
	15'h3950: q<=8'h85;
	15'h3951: q<=8'h3d;
	15'h3952: q<=8'ha5;
	15'h3953: q<=8'h05;
	15'h3954: q<=8'h10;
	15'h3955: q<=8'h16;
	15'h3956: q<=8'ha9;
	15'h3957: q<=8'h0e;
	15'h3958: q<=8'h85;
	15'h3959: q<=8'h01;
	15'h395a: q<=8'ha9;
	15'h395b: q<=8'h0a;
	15'h395c: q<=8'h85;
	15'h395d: q<=8'h00;
	15'h395e: q<=8'ha9;
	15'h395f: q<=8'h50;
	15'h3960: q<=8'hac;
	15'h3961: q<=8'h17;
	15'h3962: q<=8'h01;
	15'h3963: q<=8'hf0;
	15'h3964: q<=8'h02;
	15'h3965: q<=8'ha9;
	15'h3966: q<=8'h28;
	15'h3967: q<=8'h85;
	15'h3968: q<=8'h04;
	15'h3969: q<=8'h20;
	15'h396a: q<=8'hb2;
	15'h396b: q<=8'h92;
	15'h396c: q<=8'h20;
	15'h396d: q<=8'h48;
	15'h396e: q<=8'hca;
	15'h396f: q<=8'ha6;
	15'h3970: q<=8'h3d;
	15'h3971: q<=8'hb5;
	15'h3972: q<=8'h46;
	15'h3973: q<=8'h85;
	15'h3974: q<=8'h9f;
	15'h3975: q<=8'h20;
	15'h3976: q<=8'h25;
	15'h3977: q<=8'h90;
	15'h3978: q<=8'h4c;
	15'h3979: q<=8'h95;
	15'h397a: q<=8'hcd;
	15'h397b: q<=8'ha9;
	15'h397c: q<=8'h04;
	15'h397d: q<=8'h85;
	15'h397e: q<=8'h02;
	15'h397f: q<=8'ha9;
	15'h3980: q<=8'h00;
	15'h3981: q<=8'h85;
	15'h3982: q<=8'h01;
	15'h3983: q<=8'ha9;
	15'h3984: q<=8'h0a;
	15'h3985: q<=8'h85;
	15'h3986: q<=8'h00;
	15'h3987: q<=8'ha9;
	15'h3988: q<=8'h14;
	15'h3989: q<=8'h85;
	15'h398a: q<=8'h04;
	15'h398b: q<=8'h60;
	15'h398c: q<=8'ha6;
	15'h398d: q<=8'h3d;
	15'h398e: q<=8'hb5;
	15'h398f: q<=8'h46;
	15'h3990: q<=8'hc9;
	15'h3991: q<=8'h62;
	15'h3992: q<=8'hb0;
	15'h3993: q<=8'h04;
	15'h3994: q<=8'hf6;
	15'h3995: q<=8'h46;
	15'h3996: q<=8'he6;
	15'h3997: q<=8'h9f;
	15'h3998: q<=8'ha9;
	15'h3999: q<=8'h18;
	15'h399a: q<=8'h85;
	15'h399b: q<=8'h00;
	15'h399c: q<=8'hbd;
	15'h399d: q<=8'h02;
	15'h399e: q<=8'h01;
	15'h399f: q<=8'hf0;
	15'h39a0: q<=8'h0b;
	15'h39a1: q<=8'h20;
	15'h39a2: q<=8'hb5;
	15'h39a3: q<=8'h91;
	15'h39a4: q<=8'ha2;
	15'h39a5: q<=8'hff;
	15'h39a6: q<=8'h20;
	15'h39a7: q<=8'h6c;
	15'h39a8: q<=8'hca;
	15'h39a9: q<=8'h20;
	15'h39aa: q<=8'hb9;
	15'h39ab: q<=8'hcc;
	15'h39ac: q<=8'h4c;
	15'h39ad: q<=8'h09;
	15'h39ae: q<=8'h90;
	15'h39af: q<=8'ha9;
	15'h39b0: q<=8'h00;
	15'h39b1: q<=8'h85;
	15'h39b2: q<=8'h04;
	15'h39b3: q<=8'ha6;
	15'h39b4: q<=8'h3d;
	15'h39b5: q<=8'hd6;
	15'h39b6: q<=8'h48;
	15'h39b7: q<=8'ha5;
	15'h39b8: q<=8'h48;
	15'h39b9: q<=8'h05;
	15'h39ba: q<=8'h49;
	15'h39bb: q<=8'hd0;
	15'h39bc: q<=8'h06;
	15'h39bd: q<=8'h20;
	15'h39be: q<=8'hf1;
	15'h39bf: q<=8'hc9;
	15'h39c0: q<=8'hb8;
	15'h39c1: q<=8'h50;
	15'h39c2: q<=8'h2d;
	15'h39c3: q<=8'ha6;
	15'h39c4: q<=8'h3d;
	15'h39c5: q<=8'hb5;
	15'h39c6: q<=8'h48;
	15'h39c7: q<=8'hd0;
	15'h39c8: q<=8'h08;
	15'h39c9: q<=8'ha9;
	15'h39ca: q<=8'h0c;
	15'h39cb: q<=8'h85;
	15'h39cc: q<=8'h01;
	15'h39cd: q<=8'ha9;
	15'h39ce: q<=8'h28;
	15'h39cf: q<=8'h85;
	15'h39d0: q<=8'h04;
	15'h39d1: q<=8'ha5;
	15'h39d2: q<=8'h3e;
	15'h39d3: q<=8'hf0;
	15'h39d4: q<=8'h06;
	15'h39d5: q<=8'ha5;
	15'h39d6: q<=8'h3f;
	15'h39d7: q<=8'h49;
	15'h39d8: q<=8'h01;
	15'h39d9: q<=8'h85;
	15'h39da: q<=8'h3f;
	15'h39db: q<=8'ha6;
	15'h39dc: q<=8'h3f;
	15'h39dd: q<=8'hb5;
	15'h39de: q<=8'h48;
	15'h39df: q<=8'hf0;
	15'h39e0: q<=8'hf0;
	15'h39e1: q<=8'ha9;
	15'h39e2: q<=8'h02;
	15'h39e3: q<=8'hb4;
	15'h39e4: q<=8'h46;
	15'h39e5: q<=8'hc8;
	15'h39e6: q<=8'hd0;
	15'h39e7: q<=8'h02;
	15'h39e8: q<=8'ha9;
	15'h39e9: q<=8'h1c;
	15'h39ea: q<=8'h85;
	15'h39eb: q<=8'h02;
	15'h39ec: q<=8'ha9;
	15'h39ed: q<=8'h0a;
	15'h39ee: q<=8'h85;
	15'h39ef: q<=8'h00;
	15'h39f0: q<=8'h60;
	15'h39f1: q<=8'ha9;
	15'h39f2: q<=8'h00;
	15'h39f3: q<=8'h8d;
	15'h39f4: q<=8'h26;
	15'h39f5: q<=8'h01;
	15'h39f6: q<=8'ha6;
	15'h39f7: q<=8'h3e;
	15'h39f8: q<=8'hb5;
	15'h39f9: q<=8'h46;
	15'h39fa: q<=8'hcd;
	15'h39fb: q<=8'h26;
	15'h39fc: q<=8'h01;
	15'h39fd: q<=8'h90;
	15'h39fe: q<=8'h03;
	15'h39ff: q<=8'h8d;
	15'h3a00: q<=8'h26;
	15'h3a01: q<=8'h01;
	15'h3a02: q<=8'hca;
	15'h3a03: q<=8'h10;
	15'h3a04: q<=8'hf3;
	15'h3a05: q<=8'hac;
	15'h3a06: q<=8'h26;
	15'h3a07: q<=8'h01;
	15'h3a08: q<=8'hf0;
	15'h3a09: q<=8'h03;
	15'h3a0a: q<=8'hce;
	15'h3a0b: q<=8'h26;
	15'h3a0c: q<=8'h01;
	15'h3a0d: q<=8'ha9;
	15'h3a0e: q<=8'h14;
	15'h3a0f: q<=8'h24;
	15'h3a10: q<=8'h05;
	15'h3a11: q<=8'h10;
	15'h3a12: q<=8'h02;
	15'h3a13: q<=8'ha9;
	15'h3a14: q<=8'h10;
	15'h3a15: q<=8'h85;
	15'h3a16: q<=8'h00;
	15'h3a17: q<=8'h60;
	15'h3a18: q<=8'ha5;
	15'h3a19: q<=8'h05;
	15'h3a1a: q<=8'h29;
	15'h3a1b: q<=8'h3f;
	15'h3a1c: q<=8'h85;
	15'h3a1d: q<=8'h05;
	15'h3a1e: q<=8'ha9;
	15'h3a1f: q<=8'h00;
	15'h3a20: q<=8'h85;
	15'h3a21: q<=8'h3e;
	15'h3a22: q<=8'ha9;
	15'h3a23: q<=8'h1a;
	15'h3a24: q<=8'h85;
	15'h3a25: q<=8'h02;
	15'h3a26: q<=8'ha9;
	15'h3a27: q<=8'h0a;
	15'h3a28: q<=8'h85;
	15'h3a29: q<=8'h00;
	15'h3a2a: q<=8'ha9;
	15'h3a2b: q<=8'ha0;
	15'h3a2c: q<=8'h85;
	15'h3a2d: q<=8'h04;
	15'h3a2e: q<=8'ha9;
	15'h3a2f: q<=8'h01;
	15'h3a30: q<=8'h8d;
	15'h3a31: q<=8'h6b;
	15'h3a32: q<=8'h01;
	15'h3a33: q<=8'ha9;
	15'h3a34: q<=8'h0a;
	15'h3a35: q<=8'h85;
	15'h3a36: q<=8'h01;
	15'h3a37: q<=8'h60;
	15'h3a38: q<=8'h80;
	15'h3a39: q<=8'h40;
	15'h3a3a: q<=8'h20;
	15'h3a3b: q<=8'h10;
	15'h3a3c: q<=8'h08;
	15'h3a3d: q<=8'h04;
	15'h3a3e: q<=8'h02;
	15'h3a3f: q<=8'h01;
	15'h3a40: q<=8'h01;
	15'h3a41: q<=8'h02;
	15'h3a42: q<=8'h04;
	15'h3a43: q<=8'h08;
	15'h3a44: q<=8'h10;
	15'h3a45: q<=8'h20;
	15'h3a46: q<=8'h40;
	15'h3a47: q<=8'h80;
	15'h3a48: q<=8'ha0;
	15'h3a49: q<=8'h10;
	15'h3a4a: q<=8'had;
	15'h3a4b: q<=8'h17;
	15'h3a4c: q<=8'h01;
	15'h3a4d: q<=8'hf0;
	15'h3a4e: q<=8'h08;
	15'h3a4f: q<=8'ha5;
	15'h3a50: q<=8'h3d;
	15'h3a51: q<=8'hf0;
	15'h3a52: q<=8'h04;
	15'h3a53: q<=8'ha9;
	15'h3a54: q<=8'h04;
	15'h3a55: q<=8'ha0;
	15'h3a56: q<=8'h08;
	15'h3a57: q<=8'h45;
	15'h3a58: q<=8'ha1;
	15'h3a59: q<=8'h29;
	15'h3a5a: q<=8'h04;
	15'h3a5b: q<=8'h45;
	15'h3a5c: q<=8'ha1;
	15'h3a5d: q<=8'h85;
	15'h3a5e: q<=8'ha1;
	15'h3a5f: q<=8'h84;
	15'h3a60: q<=8'hb4;
	15'h3a61: q<=8'h60;
	15'h3a62: q<=8'ha9;
	15'h3a63: q<=8'h00;
	15'h3a64: q<=8'ha2;
	15'h3a65: q<=8'h05;
	15'h3a66: q<=8'h95;
	15'h3a67: q<=8'h40;
	15'h3a68: q<=8'hca;
	15'h3a69: q<=8'h10;
	15'h3a6a: q<=8'hfb;
	15'h3a6b: q<=8'h60;
	15'h3a6c: q<=8'hf8;
	15'h3a6d: q<=8'h24;
	15'h3a6e: q<=8'h05;
	15'h3a6f: q<=8'h10;
	15'h3a70: q<=8'h7e;
	15'h3a71: q<=8'ha4;
	15'h3a72: q<=8'h3d;
	15'h3a73: q<=8'hf0;
	15'h3a74: q<=8'h02;
	15'h3a75: q<=8'ha0;
	15'h3a76: q<=8'h03;
	15'h3a77: q<=8'he0;
	15'h3a78: q<=8'h08;
	15'h3a79: q<=8'h90;
	15'h3a7a: q<=8'h16;
	15'h3a7b: q<=8'ha5;
	15'h3a7c: q<=8'h29;
	15'h3a7d: q<=8'h18;
	15'h3a7e: q<=8'h79;
	15'h3a7f: q<=8'h40;
	15'h3a80: q<=8'h00;
	15'h3a81: q<=8'h99;
	15'h3a82: q<=8'h40;
	15'h3a83: q<=8'h00;
	15'h3a84: q<=8'ha5;
	15'h3a85: q<=8'h2a;
	15'h3a86: q<=8'h79;
	15'h3a87: q<=8'h41;
	15'h3a88: q<=8'h00;
	15'h3a89: q<=8'h99;
	15'h3a8a: q<=8'h41;
	15'h3a8b: q<=8'h00;
	15'h3a8c: q<=8'ha5;
	15'h3a8d: q<=8'h2b;
	15'h3a8e: q<=8'hb8;
	15'h3a8f: q<=8'h50;
	15'h3a90: q<=8'h15;
	15'h3a91: q<=8'hbd;
	15'h3a92: q<=8'hf1;
	15'h3a93: q<=8'hca;
	15'h3a94: q<=8'h18;
	15'h3a95: q<=8'h79;
	15'h3a96: q<=8'h40;
	15'h3a97: q<=8'h00;
	15'h3a98: q<=8'h99;
	15'h3a99: q<=8'h40;
	15'h3a9a: q<=8'h00;
	15'h3a9b: q<=8'hbd;
	15'h3a9c: q<=8'hf9;
	15'h3a9d: q<=8'hca;
	15'h3a9e: q<=8'h79;
	15'h3a9f: q<=8'h41;
	15'h3aa0: q<=8'h00;
	15'h3aa1: q<=8'h99;
	15'h3aa2: q<=8'h41;
	15'h3aa3: q<=8'h00;
	15'h3aa4: q<=8'ha9;
	15'h3aa5: q<=8'h00;
	15'h3aa6: q<=8'h08;
	15'h3aa7: q<=8'h79;
	15'h3aa8: q<=8'h42;
	15'h3aa9: q<=8'h00;
	15'h3aaa: q<=8'h99;
	15'h3aab: q<=8'h42;
	15'h3aac: q<=8'h00;
	15'h3aad: q<=8'h28;
	15'h3aae: q<=8'hf0;
	15'h3aaf: q<=8'h0b;
	15'h3ab0: q<=8'hae;
	15'h3ab1: q<=8'h56;
	15'h3ab2: q<=8'h01;
	15'h3ab3: q<=8'hf0;
	15'h3ab4: q<=8'h06;
	15'h3ab5: q<=8'he4;
	15'h3ab6: q<=8'h2b;
	15'h3ab7: q<=8'hf0;
	15'h3ab8: q<=8'h23;
	15'h3ab9: q<=8'h90;
	15'h3aba: q<=8'h21;
	15'h3abb: q<=8'h90;
	15'h3abc: q<=8'h32;
	15'h3abd: q<=8'hae;
	15'h3abe: q<=8'h56;
	15'h3abf: q<=8'h01;
	15'h3ac0: q<=8'hf0;
	15'h3ac1: q<=8'h2c;
	15'h3ac2: q<=8'he0;
	15'h3ac3: q<=8'h03;
	15'h3ac4: q<=8'h90;
	15'h3ac5: q<=8'h0b;
	15'h3ac6: q<=8'h38;
	15'h3ac7: q<=8'hed;
	15'h3ac8: q<=8'h56;
	15'h3ac9: q<=8'h01;
	15'h3aca: q<=8'hf0;
	15'h3acb: q<=8'h10;
	15'h3acc: q<=8'hb0;
	15'h3acd: q<=8'hf8;
	15'h3ace: q<=8'hb8;
	15'h3acf: q<=8'h50;
	15'h3ad0: q<=8'h1d;
	15'h3ad1: q<=8'he0;
	15'h3ad2: q<=8'h02;
	15'h3ad3: q<=8'hd0;
	15'h3ad4: q<=8'h07;
	15'h3ad5: q<=8'h29;
	15'h3ad6: q<=8'h01;
	15'h3ad7: q<=8'hf0;
	15'h3ad8: q<=8'h03;
	15'h3ad9: q<=8'hb8;
	15'h3ada: q<=8'h50;
	15'h3adb: q<=8'h12;
	15'h3adc: q<=8'ha6;
	15'h3add: q<=8'h3d;
	15'h3ade: q<=8'hb5;
	15'h3adf: q<=8'h48;
	15'h3ae0: q<=8'hc9;
	15'h3ae1: q<=8'h06;
	15'h3ae2: q<=8'hb0;
	15'h3ae3: q<=8'h0a;
	15'h3ae4: q<=8'hf6;
	15'h3ae5: q<=8'h48;
	15'h3ae6: q<=8'h20;
	15'h3ae7: q<=8'hb9;
	15'h3ae8: q<=8'hcc;
	15'h3ae9: q<=8'ha9;
	15'h3aea: q<=8'h20;
	15'h3aeb: q<=8'h8d;
	15'h3aec: q<=8'h24;
	15'h3aed: q<=8'h01;
	15'h3aee: q<=8'h38;
	15'h3aef: q<=8'hd8;
	15'h3af0: q<=8'h60;
	15'h3af1: q<=8'h00;
	15'h3af2: q<=8'h50;
	15'h3af3: q<=8'h00;
	15'h3af4: q<=8'h00;
	15'h3af5: q<=8'h50;
	15'h3af6: q<=8'h50;
	15'h3af7: q<=8'h00;
	15'h3af8: q<=8'h50;
	15'h3af9: q<=8'h00;
	15'h3afa: q<=8'h01;
	15'h3afb: q<=8'h02;
	15'h3afc: q<=8'h01;
	15'h3afd: q<=8'h00;
	15'h3afe: q<=8'h02;
	15'h3aff: q<=8'h05;
	15'h3b00: q<=8'h07;
	15'h3b01: q<=8'h00;
	15'h3b02: q<=8'h00;
	15'h3b03: q<=8'h00;
	15'h3b04: q<=8'h00;
	15'h3b05: q<=8'h00;
	15'h3b06: q<=8'h00;
	15'h3b07: q<=8'h00;
	15'h3b08: q<=8'h00;
	15'h3b09: q<=8'h35;
	15'h3b0a: q<=8'h38;
	15'h3b0b: q<=8'h00;
	15'h3b0c: q<=8'h00;
	15'h3b0d: q<=8'h00;
	15'h3b0e: q<=8'h00;
	15'h3b0f: q<=8'h00;
	15'h3b10: q<=8'h00;
	15'h3b11: q<=8'h00;
	15'h3b12: q<=8'h00;
	15'h3b13: q<=8'h47;
	15'h3b14: q<=8'h4a;
	15'h3b15: q<=8'h00;
	15'h3b16: q<=8'h00;
	15'h3b17: q<=8'h00;
	15'h3b18: q<=8'h00;
	15'h3b19: q<=8'h00;
	15'h3b1a: q<=8'h00;
	15'h3b1b: q<=8'h00;
	15'h3b1c: q<=8'h00;
	15'h3b1d: q<=8'h00;
	15'h3b1e: q<=8'h00;
	15'h3b1f: q<=8'h00;
	15'h3b20: q<=8'h00;
	15'h3b21: q<=8'h00;
	15'h3b22: q<=8'h00;
	15'h3b23: q<=8'h00;
	15'h3b24: q<=8'h00;
	15'h3b25: q<=8'h0d;
	15'h3b26: q<=8'h10;
	15'h3b27: q<=8'h00;
	15'h3b28: q<=8'h00;
	15'h3b29: q<=8'h00;
	15'h3b2a: q<=8'h00;
	15'h3b2b: q<=8'h00;
	15'h3b2c: q<=8'h00;
	15'h3b2d: q<=8'h00;
	15'h3b2e: q<=8'h00;
	15'h3b2f: q<=8'h00;
	15'h3b30: q<=8'h00;
	15'h3b31: q<=8'h00;
	15'h3b32: q<=8'h00;
	15'h3b33: q<=8'h00;
	15'h3b34: q<=8'h00;
	15'h3b35: q<=8'h00;
	15'h3b36: q<=8'h00;
	15'h3b37: q<=8'h00;
	15'h3b38: q<=8'h00;
	15'h3b39: q<=8'h00;
	15'h3b3a: q<=8'h00;
	15'h3b3b: q<=8'h65;
	15'h3b3c: q<=8'h68;
	15'h3b3d: q<=8'h00;
	15'h3b3e: q<=8'h00;
	15'h3b3f: q<=8'h00;
	15'h3b40: q<=8'h00;
	15'h3b41: q<=8'h00;
	15'h3b42: q<=8'h00;
	15'h3b43: q<=8'h00;
	15'h3b44: q<=8'h00;
	15'h3b45: q<=8'h00;
	15'h3b46: q<=8'h00;
	15'h3b47: q<=8'h21;
	15'h3b48: q<=8'h32;
	15'h3b49: q<=8'h00;
	15'h3b4a: q<=8'h00;
	15'h3b4b: q<=8'h00;
	15'h3b4c: q<=8'h00;
	15'h3b4d: q<=8'h00;
	15'h3b4e: q<=8'h00;
	15'h3b4f: q<=8'h00;
	15'h3b50: q<=8'h00;
	15'h3b51: q<=8'h13;
	15'h3b52: q<=8'h1a;
	15'h3b53: q<=8'h00;
	15'h3b54: q<=8'h00;
	15'h3b55: q<=8'h00;
	15'h3b56: q<=8'h00;
	15'h3b57: q<=8'h00;
	15'h3b58: q<=8'h00;
	15'h3b59: q<=8'h00;
	15'h3b5a: q<=8'h00;
	15'h3b5b: q<=8'h00;
	15'h3b5c: q<=8'h00;
	15'h3b5d: q<=8'h00;
	15'h3b5e: q<=8'h00;
	15'h3b5f: q<=8'h00;
	15'h3b60: q<=8'h00;
	15'h3b61: q<=8'h00;
	15'h3b62: q<=8'h00;
	15'h3b63: q<=8'h00;
	15'h3b64: q<=8'h00;
	15'h3b65: q<=8'h00;
	15'h3b66: q<=8'h00;
	15'h3b67: q<=8'h00;
	15'h3b68: q<=8'h00;
	15'h3b69: q<=8'h00;
	15'h3b6a: q<=8'h00;
	15'h3b6b: q<=8'h53;
	15'h3b6c: q<=8'h56;
	15'h3b6d: q<=8'h00;
	15'h3b6e: q<=8'h00;
	15'h3b6f: q<=8'h00;
	15'h3b70: q<=8'h00;
	15'h3b71: q<=8'h00;
	15'h3b72: q<=8'h00;
	15'h3b73: q<=8'h00;
	15'h3b74: q<=8'h00;
	15'h3b75: q<=8'h00;
	15'h3b76: q<=8'h00;
	15'h3b77: q<=8'h00;
	15'h3b78: q<=8'h00;
	15'h3b79: q<=8'h00;
	15'h3b7a: q<=8'h00;
	15'h3b7b: q<=8'h59;
	15'h3b7c: q<=8'h5c;
	15'h3b7d: q<=8'h00;
	15'h3b7e: q<=8'h00;
	15'h3b7f: q<=8'h00;
	15'h3b80: q<=8'h00;
	15'h3b81: q<=8'h00;
	15'h3b82: q<=8'h00;
	15'h3b83: q<=8'h00;
	15'h3b84: q<=8'h00;
	15'h3b85: q<=8'h00;
	15'h3b86: q<=8'h00;
	15'h3b87: q<=8'h00;
	15'h3b88: q<=8'h00;
	15'h3b89: q<=8'h00;
	15'h3b8a: q<=8'h00;
	15'h3b8b: q<=8'h00;
	15'h3b8c: q<=8'h00;
	15'h3b8d: q<=8'h00;
	15'h3b8e: q<=8'h00;
	15'h3b8f: q<=8'h3b;
	15'h3b90: q<=8'h3e;
	15'h3b91: q<=8'h00;
	15'h3b92: q<=8'h00;
	15'h3b93: q<=8'h00;
	15'h3b94: q<=8'h00;
	15'h3b95: q<=8'h00;
	15'h3b96: q<=8'h00;
	15'h3b97: q<=8'h00;
	15'h3b98: q<=8'h00;
	15'h3b99: q<=8'h00;
	15'h3b9a: q<=8'h00;
	15'h3b9b: q<=8'h00;
	15'h3b9c: q<=8'h00;
	15'h3b9d: q<=8'h41;
	15'h3b9e: q<=8'h44;
	15'h3b9f: q<=8'h00;
	15'h3ba0: q<=8'h00;
	15'h3ba1: q<=8'h4d;
	15'h3ba2: q<=8'h50;
	15'h3ba3: q<=8'h00;
	15'h3ba4: q<=8'h00;
	15'h3ba5: q<=8'h00;
	15'h3ba6: q<=8'h00;
	15'h3ba7: q<=8'h00;
	15'h3ba8: q<=8'h00;
	15'h3ba9: q<=8'h00;
	15'h3baa: q<=8'h00;
	15'h3bab: q<=8'h00;
	15'h3bac: q<=8'h00;
	15'h3bad: q<=8'h00;
	15'h3bae: q<=8'h00;
	15'h3baf: q<=8'h00;
	15'h3bb0: q<=8'h00;
	15'h3bb1: q<=8'h5f;
	15'h3bb2: q<=8'h62;
	15'h3bb3: q<=8'h00;
	15'h3bb4: q<=8'h00;
	15'h3bb5: q<=8'h00;
	15'h3bb6: q<=8'h00;
	15'h3bb7: q<=8'h00;
	15'h3bb8: q<=8'h00;
	15'h3bb9: q<=8'h00;
	15'h3bba: q<=8'h00;
	15'h3bbb: q<=8'h00;
	15'h3bbc: q<=8'h00;
	15'h3bbd: q<=8'h00;
	15'h3bbe: q<=8'h00;
	15'h3bbf: q<=8'h00;
	15'h3bc0: q<=8'h00;
	15'h3bc1: q<=8'h00;
	15'h3bc2: q<=8'h00;
	15'h3bc3: q<=8'h00;
	15'h3bc4: q<=8'h00;
	15'h3bc5: q<=8'h00;
	15'h3bc6: q<=8'h00;
	15'h3bc7: q<=8'h00;
	15'h3bc8: q<=8'h00;
	15'h3bc9: q<=8'h00;
	15'h3bca: q<=8'h00;
	15'h3bcb: q<=8'h6d;
	15'h3bcc: q<=8'h6d;
	15'h3bcd: q<=8'h00;
	15'h3bce: q<=8'h00;
	15'h3bcf: q<=8'h00;
	15'h3bd0: q<=8'h00;
	15'h3bd1: q<=8'hc0;
	15'h3bd2: q<=8'h08;
	15'h3bd3: q<=8'h04;
	15'h3bd4: q<=8'h10;
	15'h3bd5: q<=8'h00;
	15'h3bd6: q<=8'h00;
	15'h3bd7: q<=8'ha6;
	15'h3bd8: q<=8'h20;
	15'h3bd9: q<=8'hf8;
	15'h3bda: q<=8'h04;
	15'h3bdb: q<=8'h00;
	15'h3bdc: q<=8'h00;
	15'h3bdd: q<=8'h40;
	15'h3bde: q<=8'h08;
	15'h3bdf: q<=8'h04;
	15'h3be0: q<=8'h10;
	15'h3be1: q<=8'h00;
	15'h3be2: q<=8'h00;
	15'h3be3: q<=8'ha6;
	15'h3be4: q<=8'h20;
	15'h3be5: q<=8'hfe;
	15'h3be6: q<=8'h04;
	15'h3be7: q<=8'h00;
	15'h3be8: q<=8'h00;
	15'h3be9: q<=8'h10;
	15'h3bea: q<=8'h01;
	15'h3beb: q<=8'h07;
	15'h3bec: q<=8'h20;
	15'h3bed: q<=8'h00;
	15'h3bee: q<=8'h00;
	15'h3bef: q<=8'ha2;
	15'h3bf0: q<=8'h01;
	15'h3bf1: q<=8'hf8;
	15'h3bf2: q<=8'h20;
	15'h3bf3: q<=8'h00;
	15'h3bf4: q<=8'h00;
	15'h3bf5: q<=8'h08;
	15'h3bf6: q<=8'h04;
	15'h3bf7: q<=8'h20;
	15'h3bf8: q<=8'h0a;
	15'h3bf9: q<=8'h08;
	15'h3bfa: q<=8'h04;
	15'h3bfb: q<=8'h01;
	15'h3bfc: q<=8'h09;
	15'h3bfd: q<=8'h10;
	15'h3bfe: q<=8'h0d;
	15'h3bff: q<=8'h04;
	15'h3c00: q<=8'h0c;
	15'h3c01: q<=8'h00;
	15'h3c02: q<=8'h00;
	15'h3c03: q<=8'h08;
	15'h3c04: q<=8'h04;
	15'h3c05: q<=8'h00;
	15'h3c06: q<=8'h0a;
	15'h3c07: q<=8'h68;
	15'h3c08: q<=8'h04;
	15'h3c09: q<=8'h00;
	15'h3c0a: q<=8'h09;
	15'h3c0b: q<=8'h68;
	15'h3c0c: q<=8'h12;
	15'h3c0d: q<=8'hff;
	15'h3c0e: q<=8'h09;
	15'h3c0f: q<=8'h00;
	15'h3c10: q<=8'h00;
	15'h3c11: q<=8'h40;
	15'h3c12: q<=8'h01;
	15'h3c13: q<=8'h00;
	15'h3c14: q<=8'h01;
	15'h3c15: q<=8'h40;
	15'h3c16: q<=8'h01;
	15'h3c17: q<=8'hff;
	15'h3c18: q<=8'h40;
	15'h3c19: q<=8'h30;
	15'h3c1a: q<=8'h01;
	15'h3c1b: q<=8'hff;
	15'h3c1c: q<=8'h30;
	15'h3c1d: q<=8'h20;
	15'h3c1e: q<=8'h01;
	15'h3c1f: q<=8'hff;
	15'h3c20: q<=8'h20;
	15'h3c21: q<=8'h18;
	15'h3c22: q<=8'h01;
	15'h3c23: q<=8'hff;
	15'h3c24: q<=8'h18;
	15'h3c25: q<=8'h14;
	15'h3c26: q<=8'h01;
	15'h3c27: q<=8'hff;
	15'h3c28: q<=8'h14;
	15'h3c29: q<=8'h12;
	15'h3c2a: q<=8'h01;
	15'h3c2b: q<=8'hff;
	15'h3c2c: q<=8'h12;
	15'h3c2d: q<=8'h10;
	15'h3c2e: q<=8'h01;
	15'h3c2f: q<=8'hff;
	15'h3c30: q<=8'h10;
	15'h3c31: q<=8'h00;
	15'h3c32: q<=8'h00;
	15'h3c33: q<=8'ha8;
	15'h3c34: q<=8'h93;
	15'h3c35: q<=8'h00;
	15'h3c36: q<=8'h02;
	15'h3c37: q<=8'h00;
	15'h3c38: q<=8'h00;
	15'h3c39: q<=8'h0f;
	15'h3c3a: q<=8'h04;
	15'h3c3b: q<=8'h00;
	15'h3c3c: q<=8'h01;
	15'h3c3d: q<=8'h00;
	15'h3c3e: q<=8'h00;
	15'h3c3f: q<=8'ha2;
	15'h3c40: q<=8'h04;
	15'h3c41: q<=8'h40;
	15'h3c42: q<=8'h01;
	15'h3c43: q<=8'h00;
	15'h3c44: q<=8'h00;
	15'h3c45: q<=8'h00;
	15'h3c46: q<=8'h03;
	15'h3c47: q<=8'h02;
	15'h3c48: q<=8'h09;
	15'h3c49: q<=8'h00;
	15'h3c4a: q<=8'h00;
	15'h3c4b: q<=8'h08;
	15'h3c4c: q<=8'h03;
	15'h3c4d: q<=8'hff;
	15'h3c4e: q<=8'h09;
	15'h3c4f: q<=8'h00;
	15'h3c50: q<=8'h00;
	15'h3c51: q<=8'h80;
	15'h3c52: q<=8'h01;
	15'h3c53: q<=8'he8;
	15'h3c54: q<=8'h05;
	15'h3c55: q<=8'h00;
	15'h3c56: q<=8'h00;
	15'h3c57: q<=8'ha1;
	15'h3c58: q<=8'h01;
	15'h3c59: q<=8'h01;
	15'h3c5a: q<=8'h05;
	15'h3c5b: q<=8'h00;
	15'h3c5c: q<=8'h00;
	15'h3c5d: q<=8'h01;
	15'h3c5e: q<=8'h08;
	15'h3c5f: q<=8'h02;
	15'h3c60: q<=8'h10;
	15'h3c61: q<=8'h00;
	15'h3c62: q<=8'h00;
	15'h3c63: q<=8'h86;
	15'h3c64: q<=8'h20;
	15'h3c65: q<=8'h00;
	15'h3c66: q<=8'h04;
	15'h3c67: q<=8'h00;
	15'h3c68: q<=8'h00;
	15'h3c69: q<=8'h18;
	15'h3c6a: q<=8'h04;
	15'h3c6b: q<=8'h00;
	15'h3c6c: q<=8'hff;
	15'h3c6d: q<=8'h00;
	15'h3c6e: q<=8'h00;
	15'h3c6f: q<=8'haf;
	15'h3c70: q<=8'h04;
	15'h3c71: q<=8'h00;
	15'h3c72: q<=8'hff;
	15'h3c73: q<=8'h00;
	15'h3c74: q<=8'h00;
	15'h3c75: q<=8'hc0;
	15'h3c76: q<=8'h02;
	15'h3c77: q<=8'hff;
	15'h3c78: q<=8'hff;
	15'h3c79: q<=8'h00;
	15'h3c7a: q<=8'h00;
	15'h3c7b: q<=8'h28;
	15'h3c7c: q<=8'h02;
	15'h3c7d: q<=8'h00;
	15'h3c7e: q<=8'hf0;
	15'h3c7f: q<=8'h00;
	15'h3c80: q<=8'h00;
	15'h3c81: q<=8'h10;
	15'h3c82: q<=8'h0b;
	15'h3c83: q<=8'h01;
	15'h3c84: q<=8'h40;
	15'h3c85: q<=8'h00;
	15'h3c86: q<=8'h00;
	15'h3c87: q<=8'h86;
	15'h3c88: q<=8'h40;
	15'h3c89: q<=8'h00;
	15'h3c8a: q<=8'h0b;
	15'h3c8b: q<=8'h00;
	15'h3c8c: q<=8'h00;
	15'h3c8d: q<=8'h20;
	15'h3c8e: q<=8'h80;
	15'h3c8f: q<=8'h00;
	15'h3c90: q<=8'h03;
	15'h3c91: q<=8'h00;
	15'h3c92: q<=8'h00;
	15'h3c93: q<=8'ha8;
	15'h3c94: q<=8'h40;
	15'h3c95: q<=8'hf8;
	15'h3c96: q<=8'h06;
	15'h3c97: q<=8'h00;
	15'h3c98: q<=8'h00;
	15'h3c99: q<=8'hb0;
	15'h3c9a: q<=8'h02;
	15'h3c9b: q<=8'h00;
	15'h3c9c: q<=8'hff;
	15'h3c9d: q<=8'h00;
	15'h3c9e: q<=8'h00;
	15'h3c9f: q<=8'hc8;
	15'h3ca0: q<=8'h01;
	15'h3ca1: q<=8'h02;
	15'h3ca2: q<=8'hff;
	15'h3ca3: q<=8'hc8;
	15'h3ca4: q<=8'h01;
	15'h3ca5: q<=8'h02;
	15'h3ca6: q<=8'hff;
	15'h3ca7: q<=8'h00;
	15'h3ca8: q<=8'h00;
	15'h3ca9: q<=8'hc0;
	15'h3caa: q<=8'h01;
	15'h3cab: q<=8'h00;
	15'h3cac: q<=8'h01;
	15'h3cad: q<=8'h00;
	15'h3cae: q<=8'h00;
	15'h3caf: q<=8'h00;
	15'h3cb0: q<=8'ha9;
	15'h3cb1: q<=8'h5f;
	15'h3cb2: q<=8'h4c;
	15'h3cb3: q<=8'hc3;
	15'h3cb4: q<=8'hcc;
	15'h3cb5: q<=8'ha9;
	15'h3cb6: q<=8'h0f;
	15'h3cb7: q<=8'hd0;
	15'h3cb8: q<=8'h0a;
	15'h3cb9: q<=8'ha9;
	15'h3cba: q<=8'h4f;
	15'h3cbb: q<=8'hd0;
	15'h3cbc: q<=8'h06;
	15'h3cbd: q<=8'ha9;
	15'h3cbe: q<=8'h8f;
	15'h3cbf: q<=8'hd0;
	15'h3cc0: q<=8'h02;
	15'h3cc1: q<=8'ha9;
	15'h3cc2: q<=8'h1f;
	15'h3cc3: q<=8'h24;
	15'h3cc4: q<=8'h05;
	15'h3cc5: q<=8'h10;
	15'h3cc6: q<=8'h22;
	15'h3cc7: q<=8'h86;
	15'h3cc8: q<=8'h31;
	15'h3cc9: q<=8'h84;
	15'h3cca: q<=8'h32;
	15'h3ccb: q<=8'ha8;
	15'h3ccc: q<=8'ha2;
	15'h3ccd: q<=8'h0f;
	15'h3cce: q<=8'hb9;
	15'h3ccf: q<=8'h01;
	15'h3cd0: q<=8'hcb;
	15'h3cd1: q<=8'hf0;
	15'h3cd2: q<=8'h0e;
	15'h3cd3: q<=8'h86;
	15'h3cd4: q<=8'hbf;
	15'h3cd5: q<=8'h95;
	15'h3cd6: q<=8'hc0;
	15'h3cd7: q<=8'ha9;
	15'h3cd8: q<=8'h01;
	15'h3cd9: q<=8'h95;
	15'h3cda: q<=8'he0;
	15'h3cdb: q<=8'h95;
	15'h3cdc: q<=8'hf0;
	15'h3cdd: q<=8'ha9;
	15'h3cde: q<=8'hff;
	15'h3cdf: q<=8'h85;
	15'h3ce0: q<=8'hbf;
	15'h3ce1: q<=8'h88;
	15'h3ce2: q<=8'hca;
	15'h3ce3: q<=8'h10;
	15'h3ce4: q<=8'he9;
	15'h3ce5: q<=8'ha6;
	15'h3ce6: q<=8'h31;
	15'h3ce7: q<=8'ha4;
	15'h3ce8: q<=8'h32;
	15'h3ce9: q<=8'h60;
	15'h3cea: q<=8'ha9;
	15'h3ceb: q<=8'h2f;
	15'h3cec: q<=8'hd0;
	15'h3ced: q<=8'hd5;
	15'h3cee: q<=8'ha9;
	15'h3cef: q<=8'h6f;
	15'h3cf0: q<=8'hd0;
	15'h3cf1: q<=8'hd1;
	15'h3cf2: q<=8'ha9;
	15'h3cf3: q<=8'h7f;
	15'h3cf4: q<=8'hd0;
	15'h3cf5: q<=8'hcd;
	15'h3cf6: q<=8'ha9;
	15'h3cf7: q<=8'h9f;
	15'h3cf8: q<=8'hd0;
	15'h3cf9: q<=8'hc9;
	15'h3cfa: q<=8'ha9;
	15'h3cfb: q<=8'haf;
	15'h3cfc: q<=8'hd0;
	15'h3cfd: q<=8'hc9;
	15'h3cfe: q<=8'ha9;
	15'h3cff: q<=8'hbf;
	15'h3d00: q<=8'hd0;
	15'h3d01: q<=8'hc1;
	15'h3d02: q<=8'ha9;
	15'h3d03: q<=8'h3f;
	15'h3d04: q<=8'hd0;
	15'h3d05: q<=8'hbd;
	15'h3d06: q<=8'ha9;
	15'h3d07: q<=8'hcf;
	15'h3d08: q<=8'hd0;
	15'h3d09: q<=8'hb9;
	15'h3d0a: q<=8'ha2;
	15'h3d0b: q<=8'h0f;
	15'h3d0c: q<=8'hb5;
	15'h3d0d: q<=8'hc0;
	15'h3d0e: q<=8'hf0;
	15'h3d0f: q<=8'h7e;
	15'h3d10: q<=8'he4;
	15'h3d11: q<=8'hbf;
	15'h3d12: q<=8'hf0;
	15'h3d13: q<=8'h7a;
	15'h3d14: q<=8'hd6;
	15'h3d15: q<=8'he0;
	15'h3d16: q<=8'hd0;
	15'h3d17: q<=8'h76;
	15'h3d18: q<=8'hd6;
	15'h3d19: q<=8'hf0;
	15'h3d1a: q<=8'hd0;
	15'h3d1b: q<=8'h38;
	15'h3d1c: q<=8'hf6;
	15'h3d1d: q<=8'hc0;
	15'h3d1e: q<=8'hf6;
	15'h3d1f: q<=8'hc0;
	15'h3d20: q<=8'hb5;
	15'h3d21: q<=8'hc0;
	15'h3d22: q<=8'h0a;
	15'h3d23: q<=8'ha8;
	15'h3d24: q<=8'hb0;
	15'h3d25: q<=8'h10;
	15'h3d26: q<=8'hb9;
	15'h3d27: q<=8'hcb;
	15'h3d28: q<=8'hcb;
	15'h3d29: q<=8'h95;
	15'h3d2a: q<=8'hd0;
	15'h3d2b: q<=8'hb9;
	15'h3d2c: q<=8'hce;
	15'h3d2d: q<=8'hcb;
	15'h3d2e: q<=8'h95;
	15'h3d2f: q<=8'hf0;
	15'h3d30: q<=8'hb9;
	15'h3d31: q<=8'hcc;
	15'h3d32: q<=8'hcb;
	15'h3d33: q<=8'hb8;
	15'h3d34: q<=8'h50;
	15'h3d35: q<=8'h0d;
	15'h3d36: q<=8'hb9;
	15'h3d37: q<=8'hcb;
	15'h3d38: q<=8'hcc;
	15'h3d39: q<=8'h95;
	15'h3d3a: q<=8'hd0;
	15'h3d3b: q<=8'hb9;
	15'h3d3c: q<=8'hce;
	15'h3d3d: q<=8'hcc;
	15'h3d3e: q<=8'h95;
	15'h3d3f: q<=8'hf0;
	15'h3d40: q<=8'hb9;
	15'h3d41: q<=8'hcc;
	15'h3d42: q<=8'hcc;
	15'h3d43: q<=8'h95;
	15'h3d44: q<=8'he0;
	15'h3d45: q<=8'hd0;
	15'h3d46: q<=8'h0a;
	15'h3d47: q<=8'h95;
	15'h3d48: q<=8'hc0;
	15'h3d49: q<=8'hb5;
	15'h3d4a: q<=8'hd0;
	15'h3d4b: q<=8'hf0;
	15'h3d4c: q<=8'h04;
	15'h3d4d: q<=8'h95;
	15'h3d4e: q<=8'hc0;
	15'h3d4f: q<=8'hd0;
	15'h3d50: q<=8'hcb;
	15'h3d51: q<=8'hb8;
	15'h3d52: q<=8'h50;
	15'h3d53: q<=8'h2b;
	15'h3d54: q<=8'h0a;
	15'h3d55: q<=8'ha8;
	15'h3d56: q<=8'hb0;
	15'h3d57: q<=8'h0b;
	15'h3d58: q<=8'hb9;
	15'h3d59: q<=8'hcc;
	15'h3d5a: q<=8'hcb;
	15'h3d5b: q<=8'h95;
	15'h3d5c: q<=8'he0;
	15'h3d5d: q<=8'hb9;
	15'h3d5e: q<=8'hcd;
	15'h3d5f: q<=8'hcb;
	15'h3d60: q<=8'hb8;
	15'h3d61: q<=8'h50;
	15'h3d62: q<=8'h08;
	15'h3d63: q<=8'hb9;
	15'h3d64: q<=8'hcc;
	15'h3d65: q<=8'hcc;
	15'h3d66: q<=8'h95;
	15'h3d67: q<=8'he0;
	15'h3d68: q<=8'hb9;
	15'h3d69: q<=8'hcd;
	15'h3d6a: q<=8'hcc;
	15'h3d6b: q<=8'hb4;
	15'h3d6c: q<=8'hd0;
	15'h3d6d: q<=8'h18;
	15'h3d6e: q<=8'h75;
	15'h3d6f: q<=8'hd0;
	15'h3d70: q<=8'h95;
	15'h3d71: q<=8'hd0;
	15'h3d72: q<=8'h8a;
	15'h3d73: q<=8'h4a;
	15'h3d74: q<=8'h90;
	15'h3d75: q<=8'h09;
	15'h3d76: q<=8'h98;
	15'h3d77: q<=8'h55;
	15'h3d78: q<=8'hd0;
	15'h3d79: q<=8'h29;
	15'h3d7a: q<=8'hf0;
	15'h3d7b: q<=8'h55;
	15'h3d7c: q<=8'hd0;
	15'h3d7d: q<=8'h95;
	15'h3d7e: q<=8'hd0;
	15'h3d7f: q<=8'hb5;
	15'h3d80: q<=8'hd0;
	15'h3d81: q<=8'he0;
	15'h3d82: q<=8'h08;
	15'h3d83: q<=8'h90;
	15'h3d84: q<=8'h06;
	15'h3d85: q<=8'h9d;
	15'h3d86: q<=8'hc8;
	15'h3d87: q<=8'h60;
	15'h3d88: q<=8'hb8;
	15'h3d89: q<=8'h50;
	15'h3d8a: q<=8'h03;
	15'h3d8b: q<=8'h9d;
	15'h3d8c: q<=8'hc0;
	15'h3d8d: q<=8'h60;
	15'h3d8e: q<=8'hca;
	15'h3d8f: q<=8'h30;
	15'h3d90: q<=8'h03;
	15'h3d91: q<=8'h4c;
	15'h3d92: q<=8'h0c;
	15'h3d93: q<=8'hcd;
	15'h3d94: q<=8'h60;
	15'h3d95: q<=8'ha9;
	15'h3d96: q<=8'h00;
	15'h3d97: q<=8'h8d;
	15'h3d98: q<=8'hcf;
	15'h3d99: q<=8'h60;
	15'h3d9a: q<=8'h8d;
	15'h3d9b: q<=8'hdf;
	15'h3d9c: q<=8'h60;
	15'h3d9d: q<=8'h8d;
	15'h3d9e: q<=8'h20;
	15'h3d9f: q<=8'h07;
	15'h3da0: q<=8'ha2;
	15'h3da1: q<=8'h04;
	15'h3da2: q<=8'had;
	15'h3da3: q<=8'hca;
	15'h3da4: q<=8'h60;
	15'h3da5: q<=8'hac;
	15'h3da6: q<=8'hda;
	15'h3da7: q<=8'h60;
	15'h3da8: q<=8'hcd;
	15'h3da9: q<=8'hca;
	15'h3daa: q<=8'h60;
	15'h3dab: q<=8'hd0;
	15'h3dac: q<=8'h03;
	15'h3dad: q<=8'hcc;
	15'h3dae: q<=8'hda;
	15'h3daf: q<=8'h60;
	15'h3db0: q<=8'hf0;
	15'h3db1: q<=8'h05;
	15'h3db2: q<=8'h8d;
	15'h3db3: q<=8'h20;
	15'h3db4: q<=8'h07;
	15'h3db5: q<=8'ha2;
	15'h3db6: q<=8'h00;
	15'h3db7: q<=8'hca;
	15'h3db8: q<=8'h10;
	15'h3db9: q<=8'hee;
	15'h3dba: q<=8'ha9;
	15'h3dbb: q<=8'h07;
	15'h3dbc: q<=8'h8d;
	15'h3dbd: q<=8'hcf;
	15'h3dbe: q<=8'h60;
	15'h3dbf: q<=8'h8d;
	15'h3dc0: q<=8'hdf;
	15'h3dc1: q<=8'h60;
	15'h3dc2: q<=8'ha2;
	15'h3dc3: q<=8'h07;
	15'h3dc4: q<=8'ha9;
	15'h3dc5: q<=8'h00;
	15'h3dc6: q<=8'h9d;
	15'h3dc7: q<=8'hc0;
	15'h3dc8: q<=8'h60;
	15'h3dc9: q<=8'h9d;
	15'h3dca: q<=8'hd0;
	15'h3dcb: q<=8'h60;
	15'h3dcc: q<=8'h95;
	15'h3dcd: q<=8'hc0;
	15'h3dce: q<=8'h95;
	15'h3dcf: q<=8'hd0;
	15'h3dd0: q<=8'hca;
	15'h3dd1: q<=8'h10;
	15'h3dd2: q<=8'hf3;
	15'h3dd3: q<=8'ha9;
	15'h3dd4: q<=8'h00;
	15'h3dd5: q<=8'h8d;
	15'h3dd6: q<=8'hc8;
	15'h3dd7: q<=8'h60;
	15'h3dd8: q<=8'ha9;
	15'h3dd9: q<=8'h00;
	15'h3dda: q<=8'h8d;
	15'h3ddb: q<=8'hd8;
	15'h3ddc: q<=8'h60;
	15'h3ddd: q<=8'h60;
	15'h3dde: q<=8'h0b;
	15'h3ddf: q<=8'h5d;
	15'h3de0: q<=8'h22;
	15'h3de1: q<=8'h74;
	15'h3de2: q<=8'h0c;
	15'h3de3: q<=8'h5e;
	15'h3de4: q<=8'h34;
	15'h3de5: q<=8'h50;
	15'h3de6: q<=8'h00;
	15'h3de7: q<=8'h71;
	15'h3de8: q<=8'hc5;
	15'h3de9: q<=8'h68;
	15'h3dea: q<=8'h40;
	15'h3deb: q<=8'h80;
	15'h3dec: q<=8'h6c;
	15'h3ded: q<=8'h01;
	15'h3dee: q<=8'h40;
	15'h3def: q<=8'h1e;
	15'h3df0: q<=8'h00;
	15'h3df1: q<=8'h71;
	15'h3df2: q<=8'hb4;
	15'h3df3: q<=8'ha8;
	15'h3df4: q<=8'hb4;
	15'h3df5: q<=8'ha8;
	15'h3df6: q<=8'hb4;
	15'h3df7: q<=8'ha8;
	15'h3df8: q<=8'hb4;
	15'h3df9: q<=8'ha8;
	15'h3dfa: q<=8'hb4;
	15'h3dfb: q<=8'ha8;
	15'h3dfc: q<=8'h65;
	15'h3dfd: q<=8'ha8;
	15'h3dfe: q<=8'h00;
	15'h3dff: q<=8'h00;
	15'h3e00: q<=8'h70;
	15'h3e01: q<=8'h1f;
	15'h3e02: q<=8'h00;
	15'h3e03: q<=8'h71;
	15'h3e04: q<=8'h00;
	15'h3e05: q<=8'h58;
	15'h3e06: q<=8'hc1;
	15'h3e07: q<=8'h68;
	15'h3e08: q<=8'h3f;
	15'h3e09: q<=8'ha9;
	15'h3e0a: q<=8'h3f;
	15'h3e0b: q<=8'ha9;
	15'h3e0c: q<=8'h3f;
	15'h3e0d: q<=8'ha9;
	15'h3e0e: q<=8'h3f;
	15'h3e0f: q<=8'ha9;
	15'h3e10: q<=8'h3f;
	15'h3e11: q<=8'ha9;
	15'h3e12: q<=8'h3f;
	15'h3e13: q<=8'ha9;
	15'h3e14: q<=8'h30;
	15'h3e15: q<=8'h00;
	15'h3e16: q<=8'hd0;
	15'h3e17: q<=8'h1f;
	15'h3e18: q<=8'hc5;
	15'h3e19: q<=8'h68;
	15'h3e1a: q<=8'hb4;
	15'h3e1b: q<=8'ha8;
	15'h3e1c: q<=8'hb4;
	15'h3e1d: q<=8'ha8;
	15'h3e1e: q<=8'hb4;
	15'h3e1f: q<=8'ha8;
	15'h3e20: q<=8'hb4;
	15'h3e21: q<=8'ha8;
	15'h3e22: q<=8'hb4;
	15'h3e23: q<=8'ha8;
	15'h3e24: q<=8'hb4;
	15'h3e25: q<=8'ha8;
	15'h3e26: q<=8'hdc;
	15'h3e27: q<=8'h1f;
	15'h3e28: q<=8'h00;
	15'h3e29: q<=8'h00;
	15'h3e2a: q<=8'hc7;
	15'h3e2b: q<=8'h68;
	15'h3e2c: q<=8'hb4;
	15'h3e2d: q<=8'ha8;
	15'h3e2e: q<=8'hb4;
	15'h3e2f: q<=8'ha8;
	15'h3e30: q<=8'hc5;
	15'h3e31: q<=8'h68;
	15'h3e32: q<=8'h24;
	15'h3e33: q<=8'h00;
	15'h3e34: q<=8'he8;
	15'h3e35: q<=8'h1f;
	15'h3e36: q<=8'hb4;
	15'h3e37: q<=8'ha8;
	15'h3e38: q<=8'hb4;
	15'h3e39: q<=8'ha8;
	15'h3e3a: q<=8'hb4;
	15'h3e3b: q<=8'ha8;
	15'h3e3c: q<=8'h00;
	15'h3e3d: q<=8'h71;
	15'h3e3e: q<=8'he0;
	15'h3e3f: q<=8'h1f;
	15'h3e40: q<=8'h28;
	15'h3e41: q<=8'h00;
	15'h3e42: q<=8'h00;
	15'h3e43: q<=8'h71;
	15'h3e44: q<=8'hb4;
	15'h3e45: q<=8'ha8;
	15'h3e46: q<=8'hb4;
	15'h3e47: q<=8'ha8;
	15'h3e48: q<=8'hb4;
	15'h3e49: q<=8'ha8;
	15'h3e4a: q<=8'hb4;
	15'h3e4b: q<=8'ha8;
	15'h3e4c: q<=8'hb4;
	15'h3e4d: q<=8'ha8;
	15'h3e4e: q<=8'h65;
	15'h3e4f: q<=8'ha8;
	15'h3e50: q<=8'h00;
	15'h3e51: q<=8'h00;
	15'h3e52: q<=8'h70;
	15'h3e53: q<=8'h1f;
	15'h3e54: q<=8'h00;
	15'h3e55: q<=8'h71;
	15'h3e56: q<=8'h00;
	15'h3e57: q<=8'h58;
	15'h3e58: q<=8'hc1;
	15'h3e59: q<=8'h68;
	15'h3e5a: q<=8'h3f;
	15'h3e5b: q<=8'ha9;
	15'h3e5c: q<=8'h3f;
	15'h3e5d: q<=8'ha9;
	15'h3e5e: q<=8'h3f;
	15'h3e5f: q<=8'ha9;
	15'h3e60: q<=8'h3f;
	15'h3e61: q<=8'ha9;
	15'h3e62: q<=8'h3f;
	15'h3e63: q<=8'ha9;
	15'h3e64: q<=8'h3f;
	15'h3e65: q<=8'ha9;
	15'h3e66: q<=8'h55;
	15'h3e67: q<=8'h7f;
	15'h3e68: q<=8'h06;
	15'h3e69: q<=8'h20;
	15'h3e6a: q<=8'h02;
	15'h3e6b: q<=8'h22;
	15'h3e6c: q<=8'h0c;
	15'h3e6d: q<=8'h24;
	15'h3e6e: q<=8'h92;
	15'h3e6f: q<=8'h26;
	15'h3e70: q<=8'h00;
	15'h3e71: q<=8'h29;
	15'h3e72: q<=8'h56;
	15'h3e73: q<=8'h2a;
	15'h3e74: q<=8'hd8;
	15'h3e75: q<=8'h2c;
	15'h3e76: q<=8'hbe;
	15'h3e77: q<=8'h2d;
	15'h3e78: q<=8'h24;
	15'h3e79: q<=8'h2e;
	15'h3e7a: q<=8'h04;
	15'h3e7b: q<=8'h21;
	15'h3e7c: q<=8'h06;
	15'h3e7d: q<=8'h23;
	15'h3e7e: q<=8'h4e;
	15'h3e7f: q<=8'h25;
	15'h3e80: q<=8'hc8;
	15'h3e81: q<=8'h27;
	15'h3e82: q<=8'haa;
	15'h3e83: q<=8'h29;
	15'h3e84: q<=8'h96;
	15'h3e85: q<=8'h2b;
	15'h3e86: q<=8'h4a;
	15'h3e87: q<=8'h2d;
	15'h3e88: q<=8'hf0;
	15'h3e89: q<=8'h2d;
	15'h3e8a: q<=8'ha6;
	15'h3e8b: q<=8'h2e;
	15'h3e8c: q<=8'h04;
	15'h3e8d: q<=8'h20;
	15'h3e8e: q<=8'h00;
	15'h3e8f: q<=8'h22;
	15'h3e90: q<=8'h0a;
	15'h3e91: q<=8'h24;
	15'h3e92: q<=8'h90;
	15'h3e93: q<=8'h26;
	15'h3e94: q<=8'hfe;
	15'h3e95: q<=8'h28;
	15'h3e96: q<=8'h54;
	15'h3e97: q<=8'h2a;
	15'h3e98: q<=8'hd6;
	15'h3e99: q<=8'h2c;
	15'h3e9a: q<=8'hbc;
	15'h3e9b: q<=8'h2d;
	15'h3e9c: q<=8'h22;
	15'h3e9d: q<=8'h2e;
	15'h3e9e: q<=8'h03;
	15'h3e9f: q<=8'he0;
	15'h3ea0: q<=8'h01;
	15'h3ea1: q<=8'he1;
	15'h3ea2: q<=8'h06;
	15'h3ea3: q<=8'he2;
	15'h3ea4: q<=8'h49;
	15'h3ea5: q<=8'he3;
	15'h3ea6: q<=8'h80;
	15'h3ea7: q<=8'he4;
	15'h3ea8: q<=8'h2b;
	15'h3ea9: q<=8'he5;
	15'h3eaa: q<=8'h6c;
	15'h3eab: q<=8'he6;
	15'h3eac: q<=8'hdf;
	15'h3ead: q<=8'he6;
	15'h3eae: q<=8'h12;
	15'h3eaf: q<=8'he7;
	15'h3eb0: q<=8'h82;
	15'h3eb1: q<=8'he0;
	15'h3eb2: q<=8'h83;
	15'h3eb3: q<=8'he1;
	15'h3eb4: q<=8'ha7;
	15'h3eb5: q<=8'he2;
	15'h3eb6: q<=8'he4;
	15'h3eb7: q<=8'he3;
	15'h3eb8: q<=8'hd5;
	15'h3eb9: q<=8'he4;
	15'h3eba: q<=8'hcb;
	15'h3ebb: q<=8'he5;
	15'h3ebc: q<=8'ha5;
	15'h3ebd: q<=8'he6;
	15'h3ebe: q<=8'hf8;
	15'h3ebf: q<=8'he6;
	15'h3ec0: q<=8'h53;
	15'h3ec1: q<=8'he7;
	15'h3ec2: q<=8'hda;
	15'h3ec3: q<=8'hee;
	15'h3ec4: q<=8'he4;
	15'h3ec5: q<=8'hee;
	15'h3ec6: q<=8'he6;
	15'h3ec7: q<=8'hee;
	15'h3ec8: q<=8'h61;
	15'h3ec9: q<=8'haa;
	15'h3eca: q<=8'h7c;
	15'h3ecb: q<=8'haa;
	15'h3ecc: q<=8'h91;
	15'h3ecd: q<=8'haa;
	15'h3ece: q<=8'had;
	15'h3ecf: q<=8'haa;
	15'h3ed0: q<=8'hca;
	15'h3ed1: q<=8'haa;
	15'h3ed2: q<=8'h14;
	15'h3ed3: q<=8'hab;
	15'h3ed4: q<=8'h6f;
	15'h3ed5: q<=8'hab;
	15'h3ed6: q<=8'hc0;
	15'h3ed7: q<=8'hab;
	15'h3ed8: q<=8'h15;
	15'h3ed9: q<=8'hac;
	15'h3eda: q<=8'h66;
	15'h3edb: q<=8'hac;
	15'h3edc: q<=8'h7d;
	15'h3edd: q<=8'hac;
	15'h3ede: q<=8'h94;
	15'h3edf: q<=8'hac;
	15'h3ee0: q<=8'hab;
	15'h3ee1: q<=8'hac;
	15'h3ee2: q<=8'hd8;
	15'h3ee3: q<=8'hac;
	15'h3ee4: q<=8'hfa;
	15'h3ee5: q<=8'hac;
	15'h3ee6: q<=8'h0d;
	15'h3ee7: q<=8'had;
	15'h3ee8: q<=8'h20;
	15'h3ee9: q<=8'had;
	15'h3eea: q<=8'h39;
	15'h3eeb: q<=8'had;
	15'h3eec: q<=8'h51;
	15'h3eed: q<=8'had;
	15'h3eee: q<=8'h6a;
	15'h3eef: q<=8'had;
	15'h3ef0: q<=8'h8c;
	15'h3ef1: q<=8'had;
	15'h3ef2: q<=8'h8a;
	15'h3ef3: q<=8'had;
	15'h3ef4: q<=8'h88;
	15'h3ef5: q<=8'had;
	15'h3ef6: q<=8'h86;
	15'h3ef7: q<=8'had;
	15'h3ef8: q<=8'h84;
	15'h3ef9: q<=8'had;
	15'h3efa: q<=8'h82;
	15'h3efb: q<=8'had;
	15'h3efc: q<=8'h86;
	15'h3efd: q<=8'had;
	15'h3efe: q<=8'h8a;
	15'h3eff: q<=8'had;
	15'h3f00: q<=8'h8c;
	15'h3f01: q<=8'had;
	15'h3f02: q<=8'hd7;
	15'h3f03: q<=8'had;
	15'h3f04: q<=8'hc2;
	15'h3f05: q<=8'had;
	15'h3f06: q<=8'hc5;
	15'h3f07: q<=8'had;
	15'h3f08: q<=8'hc8;
	15'h3f09: q<=8'had;
	15'h3f0a: q<=8'hcb;
	15'h3f0b: q<=8'had;
	15'h3f0c: q<=8'hce;
	15'h3f0d: q<=8'had;
	15'h3f0e: q<=8'hd1;
	15'h3f0f: q<=8'had;
	15'h3f10: q<=8'hd4;
	15'h3f11: q<=8'had;
	15'h3f12: q<=8'hc2;
	15'h3f13: q<=8'hac;
	15'h3f14: q<=8'hcb;
	15'h3f15: q<=8'hac;
	15'h3f16: q<=8'h35;
	15'h3f17: q<=8'hae;
	15'h3f18: q<=8'h59;
	15'h3f19: q<=8'hae;
	15'h3f1a: q<=8'h7e;
	15'h3f1b: q<=8'hae;
	15'h3f1c: q<=8'ha2;
	15'h3f1d: q<=8'hae;
	15'h3f1e: q<=8'hc5;
	15'h3f1f: q<=8'hae;
	15'h3f20: q<=8'hcb;
	15'h3f21: q<=8'hae;
	15'h3f22: q<=8'hd2;
	15'h3f23: q<=8'hae;
	15'h3f24: q<=8'ha2;
	15'h3f25: q<=8'h02;
	15'h3f26: q<=8'had;
	15'h3f27: q<=8'h08;
	15'h3f28: q<=8'h00;
	15'h3f29: q<=8'he0;
	15'h3f2a: q<=8'h01;
	15'h3f2b: q<=8'hf0;
	15'h3f2c: q<=8'h03;
	15'h3f2d: q<=8'hb0;
	15'h3f2e: q<=8'h02;
	15'h3f2f: q<=8'h4a;
	15'h3f30: q<=8'h4a;
	15'h3f31: q<=8'h4a;
	15'h3f32: q<=8'hb5;
	15'h3f33: q<=8'h0d;
	15'h3f34: q<=8'h29;
	15'h3f35: q<=8'h1f;
	15'h3f36: q<=8'hb0;
	15'h3f37: q<=8'h37;
	15'h3f38: q<=8'hf0;
	15'h3f39: q<=8'h10;
	15'h3f3a: q<=8'hc9;
	15'h3f3b: q<=8'h1b;
	15'h3f3c: q<=8'hb0;
	15'h3f3d: q<=8'h0a;
	15'h3f3e: q<=8'ha8;
	15'h3f3f: q<=8'ha5;
	15'h3f40: q<=8'h07;
	15'h3f41: q<=8'h29;
	15'h3f42: q<=8'h07;
	15'h3f43: q<=8'hc9;
	15'h3f44: q<=8'h07;
	15'h3f45: q<=8'h98;
	15'h3f46: q<=8'h90;
	15'h3f47: q<=8'h02;
	15'h3f48: q<=8'he9;
	15'h3f49: q<=8'h01;
	15'h3f4a: q<=8'h95;
	15'h3f4b: q<=8'h0d;
	15'h3f4c: q<=8'had;
	15'h3f4d: q<=8'h08;
	15'h3f4e: q<=8'h00;
	15'h3f4f: q<=8'h29;
	15'h3f50: q<=8'h08;
	15'h3f51: q<=8'hd0;
	15'h3f52: q<=8'h04;
	15'h3f53: q<=8'ha9;
	15'h3f54: q<=8'hf0;
	15'h3f55: q<=8'h85;
	15'h3f56: q<=8'h0c;
	15'h3f57: q<=8'ha5;
	15'h3f58: q<=8'h0c;
	15'h3f59: q<=8'hf0;
	15'h3f5a: q<=8'h08;
	15'h3f5b: q<=8'hc6;
	15'h3f5c: q<=8'h0c;
	15'h3f5d: q<=8'ha9;
	15'h3f5e: q<=8'h00;
	15'h3f5f: q<=8'h95;
	15'h3f60: q<=8'h0d;
	15'h3f61: q<=8'h95;
	15'h3f62: q<=8'h10;
	15'h3f63: q<=8'h18;
	15'h3f64: q<=8'hb5;
	15'h3f65: q<=8'h10;
	15'h3f66: q<=8'hf0;
	15'h3f67: q<=8'h23;
	15'h3f68: q<=8'hd6;
	15'h3f69: q<=8'h10;
	15'h3f6a: q<=8'hd0;
	15'h3f6b: q<=8'h1f;
	15'h3f6c: q<=8'h38;
	15'h3f6d: q<=8'hb0;
	15'h3f6e: q<=8'h1c;
	15'h3f6f: q<=8'hc9;
	15'h3f70: q<=8'h1b;
	15'h3f71: q<=8'hb0;
	15'h3f72: q<=8'h09;
	15'h3f73: q<=8'hb5;
	15'h3f74: q<=8'h0d;
	15'h3f75: q<=8'h69;
	15'h3f76: q<=8'h20;
	15'h3f77: q<=8'h90;
	15'h3f78: q<=8'hd1;
	15'h3f79: q<=8'hf0;
	15'h3f7a: q<=8'h01;
	15'h3f7b: q<=8'h18;
	15'h3f7c: q<=8'ha9;
	15'h3f7d: q<=8'h1f;
	15'h3f7e: q<=8'hb0;
	15'h3f7f: q<=8'hca;
	15'h3f80: q<=8'h95;
	15'h3f81: q<=8'h0d;
	15'h3f82: q<=8'hb5;
	15'h3f83: q<=8'h10;
	15'h3f84: q<=8'hf0;
	15'h3f85: q<=8'h01;
	15'h3f86: q<=8'h38;
	15'h3f87: q<=8'ha9;
	15'h3f88: q<=8'h78;
	15'h3f89: q<=8'h95;
	15'h3f8a: q<=8'h10;
	15'h3f8b: q<=8'h90;
	15'h3f8c: q<=8'h2a;
	15'h3f8d: q<=8'ha9;
	15'h3f8e: q<=8'h00;
	15'h3f8f: q<=8'he0;
	15'h3f90: q<=8'h01;
	15'h3f91: q<=8'h90;
	15'h3f92: q<=8'h16;
	15'h3f93: q<=8'hf0;
	15'h3f94: q<=8'h0c;
	15'h3f95: q<=8'ha5;
	15'h3f96: q<=8'h09;
	15'h3f97: q<=8'h29;
	15'h3f98: q<=8'h0c;
	15'h3f99: q<=8'h4a;
	15'h3f9a: q<=8'h4a;
	15'h3f9b: q<=8'hf0;
	15'h3f9c: q<=8'h0c;
	15'h3f9d: q<=8'h69;
	15'h3f9e: q<=8'h02;
	15'h3f9f: q<=8'hd0;
	15'h3fa0: q<=8'h08;
	15'h3fa1: q<=8'ha5;
	15'h3fa2: q<=8'h09;
	15'h3fa3: q<=8'h29;
	15'h3fa4: q<=8'h10;
	15'h3fa5: q<=8'hf0;
	15'h3fa6: q<=8'h02;
	15'h3fa7: q<=8'ha9;
	15'h3fa8: q<=8'h01;
	15'h3fa9: q<=8'h38;
	15'h3faa: q<=8'h48;
	15'h3fab: q<=8'h65;
	15'h3fac: q<=8'h16;
	15'h3fad: q<=8'h85;
	15'h3fae: q<=8'h16;
	15'h3faf: q<=8'h68;
	15'h3fb0: q<=8'h38;
	15'h3fb1: q<=8'h65;
	15'h3fb2: q<=8'h17;
	15'h3fb3: q<=8'h85;
	15'h3fb4: q<=8'h17;
	15'h3fb5: q<=8'hf6;
	15'h3fb6: q<=8'h13;
	15'h3fb7: q<=8'hca;
	15'h3fb8: q<=8'h30;
	15'h3fb9: q<=8'h03;
	15'h3fba: q<=8'h4c;
	15'h3fbb: q<=8'h26;
	15'h3fbc: q<=8'hcf;
	15'h3fbd: q<=8'ha5;
	15'h3fbe: q<=8'h09;
	15'h3fbf: q<=8'h4a;
	15'h3fc0: q<=8'h4a;
	15'h3fc1: q<=8'h4a;
	15'h3fc2: q<=8'h4a;
	15'h3fc3: q<=8'h4a;
	15'h3fc4: q<=8'ha8;
	15'h3fc5: q<=8'ha5;
	15'h3fc6: q<=8'h16;
	15'h3fc7: q<=8'h38;
	15'h3fc8: q<=8'hf9;
	15'h3fc9: q<=8'hd9;
	15'h3fca: q<=8'hcf;
	15'h3fcb: q<=8'h30;
	15'h3fcc: q<=8'h14;
	15'h3fcd: q<=8'h85;
	15'h3fce: q<=8'h16;
	15'h3fcf: q<=8'he6;
	15'h3fd0: q<=8'h18;
	15'h3fd1: q<=8'hc0;
	15'h3fd2: q<=8'h03;
	15'h3fd3: q<=8'hd0;
	15'h3fd4: q<=8'h0c;
	15'h3fd5: q<=8'he6;
	15'h3fd6: q<=8'h18;
	15'h3fd7: q<=8'hd0;
	15'h3fd8: q<=8'h08;
	15'h3fd9: q<=8'h7f;
	15'h3fda: q<=8'h02;
	15'h3fdb: q<=8'h04;
	15'h3fdc: q<=8'h04;
	15'h3fdd: q<=8'h05;
	15'h3fde: q<=8'h03;
	15'h3fdf: q<=8'h7f;
	15'h3fe0: q<=8'h7f;
	15'h3fe1: q<=8'ha5;
	15'h3fe2: q<=8'h09;
	15'h3fe3: q<=8'h29;
	15'h3fe4: q<=8'h03;
	15'h3fe5: q<=8'ha8;
	15'h3fe6: q<=8'hf0;
	15'h3fe7: q<=8'h1a;
	15'h3fe8: q<=8'h4a;
	15'h3fe9: q<=8'h69;
	15'h3fea: q<=8'h00;
	15'h3feb: q<=8'h49;
	15'h3fec: q<=8'hff;
	15'h3fed: q<=8'h38;
	15'h3fee: q<=8'h65;
	15'h3fef: q<=8'h17;
	15'h3ff0: q<=8'hb0;
	15'h3ff1: q<=8'h08;
	15'h3ff2: q<=8'h65;
	15'h3ff3: q<=8'h18;
	15'h3ff4: q<=8'h30;
	15'h3ff5: q<=8'h0e;
	15'h3ff6: q<=8'h85;
	15'h3ff7: q<=8'h18;
	15'h3ff8: q<=8'ha9;
	15'h3ff9: q<=8'h00;
	15'h3ffa: q<=8'hc0;
	15'h3ffb: q<=8'h02;
	15'h3ffc: q<=8'hb0;
	15'h3ffd: q<=8'h02;
	15'h3ffe: q<=8'he6;
	15'h3fff: q<=8'h06;
	15'h4000: q<=8'he6;
	15'h4001: q<=8'h06;
	15'h4002: q<=8'h85;
	15'h4003: q<=8'h17;
	15'h4004: q<=8'ha5;
	15'h4005: q<=8'h07;
	15'h4006: q<=8'h4a;
	15'h4007: q<=8'hb0;
	15'h4008: q<=8'h27;
	15'h4009: q<=8'ha0;
	15'h400a: q<=8'h00;
	15'h400b: q<=8'ha2;
	15'h400c: q<=8'h02;
	15'h400d: q<=8'hb5;
	15'h400e: q<=8'h13;
	15'h400f: q<=8'hf0;
	15'h4010: q<=8'h09;
	15'h4011: q<=8'hc9;
	15'h4012: q<=8'h10;
	15'h4013: q<=8'h90;
	15'h4014: q<=8'h05;
	15'h4015: q<=8'h69;
	15'h4016: q<=8'hef;
	15'h4017: q<=8'hc8;
	15'h4018: q<=8'h95;
	15'h4019: q<=8'h13;
	15'h401a: q<=8'hca;
	15'h401b: q<=8'h10;
	15'h401c: q<=8'hf0;
	15'h401d: q<=8'h98;
	15'h401e: q<=8'hd0;
	15'h401f: q<=8'h10;
	15'h4020: q<=8'ha2;
	15'h4021: q<=8'h02;
	15'h4022: q<=8'hb5;
	15'h4023: q<=8'h13;
	15'h4024: q<=8'hf0;
	15'h4025: q<=8'h07;
	15'h4026: q<=8'h18;
	15'h4027: q<=8'h69;
	15'h4028: q<=8'hef;
	15'h4029: q<=8'h95;
	15'h402a: q<=8'h13;
	15'h402b: q<=8'h30;
	15'h402c: q<=8'h03;
	15'h402d: q<=8'hca;
	15'h402e: q<=8'h10;
	15'h402f: q<=8'hf2;
	15'h4030: q<=8'h60;
	15'h4031: q<=8'h5d;
	15'h4032: q<=8'hd1;
	15'h4033: q<=8'h8f;
	15'h4034: q<=8'hd1;
	15'h4035: q<=8'h8f;
	15'h4036: q<=8'hd1;
	15'h4037: q<=8'hb1;
	15'h4038: q<=8'hd1;
	15'h4039: q<=8'heb;
	15'h403a: q<=8'hd1;
	15'h403b: q<=8'h03;
	15'h403c: q<=8'hd2;
	15'h403d: q<=8'h61;
	15'h403e: q<=8'hd2;
	15'h403f: q<=8'hcb;
	15'h4040: q<=8'hd2;
	15'h4041: q<=8'h33;
	15'h4042: q<=8'hd3;
	15'h4043: q<=8'h66;
	15'h4044: q<=8'hd3;
	15'h4045: q<=8'hb0;
	15'h4046: q<=8'hd3;
	15'h4047: q<=8'he6;
	15'h4048: q<=8'hd3;
	15'h4049: q<=8'hff;
	15'h404a: q<=8'hd3;
	15'h404b: q<=8'h17;
	15'h404c: q<=8'hd4;
	15'h404d: q<=8'h1d;
	15'h404e: q<=8'hd4;
	15'h404f: q<=8'h34;
	15'h4050: q<=8'hd4;
	15'h4051: q<=8'h4c;
	15'h4052: q<=8'hd4;
	15'h4053: q<=8'h60;
	15'h4054: q<=8'hd4;
	15'h4055: q<=8'ha1;
	15'h4056: q<=8'hd4;
	15'h4057: q<=8'hab;
	15'h4058: q<=8'hd4;
	15'h4059: q<=8'hef;
	15'h405a: q<=8'hd4;
	15'h405b: q<=8'h30;
	15'h405c: q<=8'hd5;
	15'h405d: q<=8'h75;
	15'h405e: q<=8'hd5;
	15'h405f: q<=8'h85;
	15'h4060: q<=8'hd5;
	15'h4061: q<=8'ha1;
	15'h4062: q<=8'hd5;
	15'h4063: q<=8'ha8;
	15'h4064: q<=8'hd5;
	15'h4065: q<=8'he9;
	15'h4066: q<=8'hd5;
	15'h4067: q<=8'h1c;
	15'h4068: q<=8'hd6;
	15'h4069: q<=8'h62;
	15'h406a: q<=8'hd6;
	15'h406b: q<=8'h7a;
	15'h406c: q<=8'hd6;
	15'h406d: q<=8'h67;
	15'h406e: q<=8'hd1;
	15'h406f: q<=8'h97;
	15'h4070: q<=8'hd1;
	15'h4071: q<=8'h97;
	15'h4072: q<=8'hd1;
	15'h4073: q<=8'hbd;
	15'h4074: q<=8'hd1;
	15'h4075: q<=8'hf0;
	15'h4076: q<=8'hd1;
	15'h4077: q<=8'h17;
	15'h4078: q<=8'hd2;
	15'h4079: q<=8'h75;
	15'h407a: q<=8'hd2;
	15'h407b: q<=8'he0;
	15'h407c: q<=8'hd2;
	15'h407d: q<=8'h3f;
	15'h407e: q<=8'hd3;
	15'h407f: q<=8'h79;
	15'h4080: q<=8'hd3;
	15'h4081: q<=8'hbe;
	15'h4082: q<=8'hd3;
	15'h4083: q<=8'he6;
	15'h4084: q<=8'hd3;
	15'h4085: q<=8'hff;
	15'h4086: q<=8'hd3;
	15'h4087: q<=8'h17;
	15'h4088: q<=8'hd4;
	15'h4089: q<=8'h22;
	15'h408a: q<=8'hd4;
	15'h408b: q<=8'h3a;
	15'h408c: q<=8'hd4;
	15'h408d: q<=8'h51;
	15'h408e: q<=8'hd4;
	15'h408f: q<=8'h6d;
	15'h4090: q<=8'hd4;
	15'h4091: q<=8'ha1;
	15'h4092: q<=8'hd4;
	15'h4093: q<=8'hba;
	15'h4094: q<=8'hd4;
	15'h4095: q<=8'hfd;
	15'h4096: q<=8'hd4;
	15'h4097: q<=8'h3f;
	15'h4098: q<=8'hd5;
	15'h4099: q<=8'h75;
	15'h409a: q<=8'hd5;
	15'h409b: q<=8'h85;
	15'h409c: q<=8'hd5;
	15'h409d: q<=8'ha1;
	15'h409e: q<=8'hd5;
	15'h409f: q<=8'hb9;
	15'h40a0: q<=8'hd5;
	15'h40a1: q<=8'hf6;
	15'h40a2: q<=8'hd5;
	15'h40a3: q<=8'h29;
	15'h40a4: q<=8'hd6;
	15'h40a5: q<=8'h68;
	15'h40a6: q<=8'hd6;
	15'h40a7: q<=8'h7a;
	15'h40a8: q<=8'hd6;
	15'h40a9: q<=8'h75;
	15'h40aa: q<=8'hd1;
	15'h40ab: q<=8'h9f;
	15'h40ac: q<=8'hd1;
	15'h40ad: q<=8'h9f;
	15'h40ae: q<=8'hd1;
	15'h40af: q<=8'hcf;
	15'h40b0: q<=8'hd1;
	15'h40b1: q<=8'hf6;
	15'h40b2: q<=8'hd1;
	15'h40b3: q<=8'h30;
	15'h40b4: q<=8'hd2;
	15'h40b5: q<=8'h94;
	15'h40b6: q<=8'hd2;
	15'h40b7: q<=8'hfb;
	15'h40b8: q<=8'hd2;
	15'h40b9: q<=8'h50;
	15'h40ba: q<=8'hd3;
	15'h40bb: q<=8'h8b;
	15'h40bc: q<=8'hd3;
	15'h40bd: q<=8'hcb;
	15'h40be: q<=8'hd3;
	15'h40bf: q<=8'hf5;
	15'h40c0: q<=8'hd3;
	15'h40c1: q<=8'h0e;
	15'h40c2: q<=8'hd4;
	15'h40c3: q<=8'h17;
	15'h40c4: q<=8'hd4;
	15'h40c5: q<=8'h28;
	15'h40c6: q<=8'hd4;
	15'h40c7: q<=8'h41;
	15'h40c8: q<=8'hd4;
	15'h40c9: q<=8'h5b;
	15'h40ca: q<=8'hd4;
	15'h40cb: q<=8'h83;
	15'h40cc: q<=8'hd4;
	15'h40cd: q<=8'ha1;
	15'h40ce: q<=8'hd4;
	15'h40cf: q<=8'hcc;
	15'h40d0: q<=8'hd4;
	15'h40d1: q<=8'h0e;
	15'h40d2: q<=8'hd5;
	15'h40d3: q<=8'h51;
	15'h40d4: q<=8'hd5;
	15'h40d5: q<=8'h75;
	15'h40d6: q<=8'hd5;
	15'h40d7: q<=8'h8e;
	15'h40d8: q<=8'hd5;
	15'h40d9: q<=8'ha1;
	15'h40da: q<=8'hd5;
	15'h40db: q<=8'hc8;
	15'h40dc: q<=8'hd5;
	15'h40dd: q<=8'h04;
	15'h40de: q<=8'hd6;
	15'h40df: q<=8'h3e;
	15'h40e0: q<=8'hd6;
	15'h40e1: q<=8'h6f;
	15'h40e2: q<=8'hd6;
	15'h40e3: q<=8'h8f;
	15'h40e4: q<=8'hd6;
	15'h40e5: q<=8'h7f;
	15'h40e6: q<=8'hd1;
	15'h40e7: q<=8'ha8;
	15'h40e8: q<=8'hd1;
	15'h40e9: q<=8'ha8;
	15'h40ea: q<=8'hd1;
	15'h40eb: q<=8'hde;
	15'h40ec: q<=8'hd1;
	15'h40ed: q<=8'hfc;
	15'h40ee: q<=8'hd1;
	15'h40ef: q<=8'h4d;
	15'h40f0: q<=8'hd2;
	15'h40f1: q<=8'hae;
	15'h40f2: q<=8'hd2;
	15'h40f3: q<=8'h16;
	15'h40f4: q<=8'hd3;
	15'h40f5: q<=8'h5e;
	15'h40f6: q<=8'hd3;
	15'h40f7: q<=8'ha0;
	15'h40f8: q<=8'hd3;
	15'h40f9: q<=8'hda;
	15'h40fa: q<=8'hd3;
	15'h40fb: q<=8'hed;
	15'h40fc: q<=8'hd3;
	15'h40fd: q<=8'h06;
	15'h40fe: q<=8'hd4;
	15'h40ff: q<=8'h17;
	15'h4100: q<=8'hd4;
	15'h4101: q<=8'h2d;
	15'h4102: q<=8'hd4;
	15'h4103: q<=8'h46;
	15'h4104: q<=8'hd4;
	15'h4105: q<=8'h56;
	15'h4106: q<=8'hd4;
	15'h4107: q<=8'h92;
	15'h4108: q<=8'hd4;
	15'h4109: q<=8'ha1;
	15'h410a: q<=8'hd4;
	15'h410b: q<=8'hdd;
	15'h410c: q<=8'hd4;
	15'h410d: q<=8'h1f;
	15'h410e: q<=8'hd5;
	15'h410f: q<=8'h63;
	15'h4110: q<=8'hd5;
	15'h4111: q<=8'h75;
	15'h4112: q<=8'hd5;
	15'h4113: q<=8'h97;
	15'h4114: q<=8'hd5;
	15'h4115: q<=8'ha1;
	15'h4116: q<=8'hd5;
	15'h4117: q<=8'hd9;
	15'h4118: q<=8'hd5;
	15'h4119: q<=8'h10;
	15'h411a: q<=8'hd6;
	15'h411b: q<=8'h51;
	15'h411c: q<=8'hd6;
	15'h411d: q<=8'h74;
	15'h411e: q<=8'hd6;
	15'h411f: q<=8'ha1;
	15'h4120: q<=8'hd6;
	15'h4121: q<=8'h51;
	15'h4122: q<=8'h56;
	15'h4123: q<=8'h00;
	15'h4124: q<=8'h1a;
	15'h4125: q<=8'h01;
	15'h4126: q<=8'h20;
	15'h4127: q<=8'h31;
	15'h4128: q<=8'h56;
	15'h4129: q<=8'h01;
	15'h412a: q<=8'h38;
	15'h412b: q<=8'h31;
	15'h412c: q<=8'hb0;
	15'h412d: q<=8'h41;
	15'h412e: q<=8'h00;
	15'h412f: q<=8'h11;
	15'h4130: q<=8'hf6;
	15'h4131: q<=8'h30;
	15'h4132: q<=8'h38;
	15'h4133: q<=8'h31;
	15'h4134: q<=8'hce;
	15'h4135: q<=8'h51;
	15'h4136: q<=8'h0a;
	15'h4137: q<=8'h31;
	15'h4138: q<=8'he2;
	15'h4139: q<=8'h31;
	15'h413a: q<=8'he2;
	15'h413b: q<=8'h51;
	15'h413c: q<=8'hba;
	15'h413d: q<=8'h51;
	15'h413e: q<=8'h98;
	15'h413f: q<=8'h51;
	15'h4140: q<=8'hd8;
	15'h4141: q<=8'h51;
	15'h4142: q<=8'hc9;
	15'h4143: q<=8'h31;
	15'h4144: q<=8'h56;
	15'h4145: q<=8'h51;
	15'h4146: q<=8'h80;
	15'h4147: q<=8'h51;
	15'h4148: q<=8'h80;
	15'h4149: q<=8'h51;
	15'h414a: q<=8'h80;
	15'h414b: q<=8'h51;
	15'h414c: q<=8'h80;
	15'h414d: q<=8'h71;
	15'h414e: q<=8'h92;
	15'h414f: q<=8'h51;
	15'h4150: q<=8'h80;
	15'h4151: q<=8'h31;
	15'h4152: q<=8'hb0;
	15'h4153: q<=8'h51;
	15'h4154: q<=8'h89;
	15'h4155: q<=8'h41;
	15'h4156: q<=8'h89;
	15'h4157: q<=8'h00;
	15'h4158: q<=8'h00;
	15'h4159: q<=8'h71;
	15'h415a: q<=8'h5a;
	15'h415b: q<=8'h71;
	15'h415c: q<=8'ha0;
	15'h415d: q<=8'he5;
	15'h415e: q<=8'h22;
	15'h415f: q<=8'h16;
	15'h4160: q<=8'h2e;
	15'h4161: q<=8'h1e;
	15'h4162: q<=8'h00;
	15'h4163: q<=8'h32;
	15'h4164: q<=8'h40;
	15'h4165: q<=8'h1e;
	15'h4166: q<=8'hb8;
	15'h4167: q<=8'hd9;
	15'h4168: q<=8'h20;
	15'h4169: q<=8'h26;
	15'h416a: q<=8'h30;
	15'h416b: q<=8'h00;
	15'h416c: q<=8'h1c;
	15'h416d: q<=8'h1e;
	15'h416e: q<=8'h00;
	15'h416f: q<=8'h34;
	15'h4170: q<=8'h16;
	15'h4171: q<=8'h38;
	15'h4172: q<=8'h3c;
	15'h4173: q<=8'h26;
	15'h4174: q<=8'h9e;
	15'h4175: q<=8'he5;
	15'h4176: q<=8'h3a;
	15'h4177: q<=8'h34;
	15'h4178: q<=8'h26;
	15'h4179: q<=8'h1e;
	15'h417a: q<=8'h2c;
	15'h417b: q<=8'h1e;
	15'h417c: q<=8'h30;
	15'h417d: q<=8'h1c;
	15'h417e: q<=8'h9e;
	15'h417f: q<=8'hd3;
	15'h4180: q<=8'h28;
	15'h4181: q<=8'h3e;
	15'h4182: q<=8'h1e;
	15'h4183: q<=8'h22;
	15'h4184: q<=8'h32;
	15'h4185: q<=8'h00;
	15'h4186: q<=8'h3c;
	15'h4187: q<=8'h1e;
	15'h4188: q<=8'h38;
	15'h4189: q<=8'h2e;
	15'h418a: q<=8'h26;
	15'h418b: q<=8'h30;
	15'h418c: q<=8'h16;
	15'h418d: q<=8'h1c;
	15'h418e: q<=8'hb2;
	15'h418f: q<=8'hcd;
	15'h4190: q<=8'h34;
	15'h4191: q<=8'h2c;
	15'h4192: q<=8'h16;
	15'h4193: q<=8'h46;
	15'h4194: q<=8'h1e;
	15'h4195: q<=8'h38;
	15'h4196: q<=8'h80;
	15'h4197: q<=8'hc6;
	15'h4198: q<=8'h28;
	15'h4199: q<=8'h32;
	15'h419a: q<=8'h3e;
	15'h419b: q<=8'h1e;
	15'h419c: q<=8'h3e;
	15'h419d: q<=8'h38;
	15'h419e: q<=8'h80;
	15'h419f: q<=8'hc6;
	15'h41a0: q<=8'h3a;
	15'h41a1: q<=8'h34;
	15'h41a2: q<=8'h26;
	15'h41a3: q<=8'h1e;
	15'h41a4: q<=8'h2c;
	15'h41a5: q<=8'h1e;
	15'h41a6: q<=8'h38;
	15'h41a7: q<=8'h80;
	15'h41a8: q<=8'hc6;
	15'h41a9: q<=8'h28;
	15'h41aa: q<=8'h3e;
	15'h41ab: q<=8'h22;
	15'h41ac: q<=8'h16;
	15'h41ad: q<=8'h1c;
	15'h41ae: q<=8'h32;
	15'h41af: q<=8'h38;
	15'h41b0: q<=8'h80;
	15'h41b1: q<=8'hdf;
	15'h41b2: q<=8'h34;
	15'h41b3: q<=8'h38;
	15'h41b4: q<=8'h1e;
	15'h41b5: q<=8'h3a;
	15'h41b6: q<=8'h3a;
	15'h41b7: q<=8'h00;
	15'h41b8: q<=8'h3a;
	15'h41b9: q<=8'h3c;
	15'h41ba: q<=8'h16;
	15'h41bb: q<=8'h38;
	15'h41bc: q<=8'hbc;
	15'h41bd: q<=8'hcd;
	15'h41be: q<=8'h16;
	15'h41bf: q<=8'h34;
	15'h41c0: q<=8'h34;
	15'h41c1: q<=8'h3e;
	15'h41c2: q<=8'h46;
	15'h41c3: q<=8'h1e;
	15'h41c4: q<=8'h48;
	15'h41c5: q<=8'h00;
	15'h41c6: q<=8'h3a;
	15'h41c7: q<=8'h3e;
	15'h41c8: q<=8'h38;
	15'h41c9: q<=8'h00;
	15'h41ca: q<=8'h3a;
	15'h41cb: q<=8'h3c;
	15'h41cc: q<=8'h16;
	15'h41cd: q<=8'h38;
	15'h41ce: q<=8'hbc;
	15'h41cf: q<=8'hd6;
	15'h41d0: q<=8'h3a;
	15'h41d1: q<=8'h3c;
	15'h41d2: q<=8'h16;
	15'h41d3: q<=8'h38;
	15'h41d4: q<=8'h3c;
	15'h41d5: q<=8'h00;
	15'h41d6: q<=8'h1c;
	15'h41d7: q<=8'h38;
	15'h41d8: q<=8'h3e;
	15'h41d9: q<=8'h1e;
	15'h41da: q<=8'h1a;
	15'h41db: q<=8'h2a;
	15'h41dc: q<=8'h1e;
	15'h41dd: q<=8'hb0;
	15'h41de: q<=8'hdc;
	15'h41df: q<=8'h34;
	15'h41e0: q<=8'h3e;
	15'h41e1: q<=8'h2c;
	15'h41e2: q<=8'h3a;
	15'h41e3: q<=8'h16;
	15'h41e4: q<=8'h38;
	15'h41e5: q<=8'h00;
	15'h41e6: q<=8'h3a;
	15'h41e7: q<=8'h3c;
	15'h41e8: q<=8'h16;
	15'h41e9: q<=8'h38;
	15'h41ea: q<=8'hbc;
	15'h41eb: q<=8'hf4;
	15'h41ec: q<=8'h34;
	15'h41ed: q<=8'h2c;
	15'h41ee: q<=8'h16;
	15'h41ef: q<=8'hc6;
	15'h41f0: q<=8'hf1;
	15'h41f1: q<=8'h28;
	15'h41f2: q<=8'h32;
	15'h41f3: q<=8'h3e;
	15'h41f4: q<=8'h1e;
	15'h41f5: q<=8'hc8;
	15'h41f6: q<=8'hf1;
	15'h41f7: q<=8'h3a;
	15'h41f8: q<=8'h34;
	15'h41f9: q<=8'h26;
	15'h41fa: q<=8'h1e;
	15'h41fb: q<=8'hac;
	15'h41fc: q<=8'hee;
	15'h41fd: q<=8'h28;
	15'h41fe: q<=8'h3e;
	15'h41ff: q<=8'h1e;
	15'h4200: q<=8'h22;
	15'h4201: q<=8'h3e;
	15'h4202: q<=8'h9e;
	15'h4203: q<=8'hc7;
	15'h4204: q<=8'h1e;
	15'h4205: q<=8'h30;
	15'h4206: q<=8'h3c;
	15'h4207: q<=8'h1e;
	15'h4208: q<=8'h38;
	15'h4209: q<=8'h00;
	15'h420a: q<=8'h46;
	15'h420b: q<=8'h32;
	15'h420c: q<=8'h3e;
	15'h420d: q<=8'h38;
	15'h420e: q<=8'h00;
	15'h420f: q<=8'h26;
	15'h4210: q<=8'h30;
	15'h4211: q<=8'h26;
	15'h4212: q<=8'h3c;
	15'h4213: q<=8'h26;
	15'h4214: q<=8'h16;
	15'h4215: q<=8'h2c;
	15'h4216: q<=8'hba;
	15'h4217: q<=8'hb8;
	15'h4218: q<=8'h3a;
	15'h4219: q<=8'h40;
	15'h421a: q<=8'h34;
	15'h421b: q<=8'h00;
	15'h421c: q<=8'h1e;
	15'h421d: q<=8'h30;
	15'h421e: q<=8'h3c;
	15'h421f: q<=8'h38;
	15'h4220: q<=8'h1e;
	15'h4221: q<=8'h48;
	15'h4222: q<=8'h00;
	15'h4223: q<=8'h40;
	15'h4224: q<=8'h32;
	15'h4225: q<=8'h3a;
	15'h4226: q<=8'h00;
	15'h4227: q<=8'h26;
	15'h4228: q<=8'h30;
	15'h4229: q<=8'h26;
	15'h422a: q<=8'h3c;
	15'h422b: q<=8'h26;
	15'h422c: q<=8'h16;
	15'h422d: q<=8'h2c;
	15'h422e: q<=8'h1e;
	15'h422f: q<=8'hba;
	15'h4230: q<=8'hac;
	15'h4231: q<=8'h22;
	15'h4232: q<=8'h1e;
	15'h4233: q<=8'h18;
	15'h4234: q<=8'h1e;
	15'h4235: q<=8'h30;
	15'h4236: q<=8'h00;
	15'h4237: q<=8'h3a;
	15'h4238: q<=8'h26;
	15'h4239: q<=8'h1e;
	15'h423a: q<=8'h00;
	15'h423b: q<=8'h26;
	15'h423c: q<=8'h24;
	15'h423d: q<=8'h38;
	15'h423e: q<=8'h1e;
	15'h423f: q<=8'h00;
	15'h4240: q<=8'h26;
	15'h4241: q<=8'h30;
	15'h4242: q<=8'h26;
	15'h4243: q<=8'h3c;
	15'h4244: q<=8'h26;
	15'h4245: q<=8'h16;
	15'h4246: q<=8'h2c;
	15'h4247: q<=8'h1e;
	15'h4248: q<=8'h30;
	15'h4249: q<=8'h00;
	15'h424a: q<=8'h1e;
	15'h424b: q<=8'h26;
	15'h424c: q<=8'hb0;
	15'h424d: q<=8'hc7;
	15'h424e: q<=8'h1e;
	15'h424f: q<=8'h30;
	15'h4250: q<=8'h3c;
	15'h4251: q<=8'h38;
	15'h4252: q<=8'h1e;
	15'h4253: q<=8'h00;
	15'h4254: q<=8'h3a;
	15'h4255: q<=8'h3e;
	15'h4256: q<=8'h3a;
	15'h4257: q<=8'h00;
	15'h4258: q<=8'h26;
	15'h4259: q<=8'h30;
	15'h425a: q<=8'h26;
	15'h425b: q<=8'h1a;
	15'h425c: q<=8'h26;
	15'h425d: q<=8'h16;
	15'h425e: q<=8'h2c;
	15'h425f: q<=8'h1e;
	15'h4260: q<=8'hba;
	15'h4261: q<=8'hc7;
	15'h4262: q<=8'h3a;
	15'h4263: q<=8'h34;
	15'h4264: q<=8'h26;
	15'h4265: q<=8'h30;
	15'h4266: q<=8'h00;
	15'h4267: q<=8'h2a;
	15'h4268: q<=8'h30;
	15'h4269: q<=8'h32;
	15'h426a: q<=8'h18;
	15'h426b: q<=8'h00;
	15'h426c: q<=8'h3c;
	15'h426d: q<=8'h32;
	15'h426e: q<=8'h00;
	15'h426f: q<=8'h1a;
	15'h4270: q<=8'h24;
	15'h4271: q<=8'h16;
	15'h4272: q<=8'h30;
	15'h4273: q<=8'h22;
	15'h4274: q<=8'h9e;
	15'h4275: q<=8'ha6;
	15'h4276: q<=8'h3c;
	15'h4277: q<=8'h32;
	15'h4278: q<=8'h3e;
	15'h4279: q<=8'h38;
	15'h427a: q<=8'h30;
	15'h427b: q<=8'h1e;
	15'h427c: q<=8'h48;
	15'h427d: q<=8'h00;
	15'h427e: q<=8'h2c;
	15'h427f: q<=8'h1e;
	15'h4280: q<=8'h00;
	15'h4281: q<=8'h18;
	15'h4282: q<=8'h32;
	15'h4283: q<=8'h3e;
	15'h4284: q<=8'h3c;
	15'h4285: q<=8'h32;
	15'h4286: q<=8'h30;
	15'h4287: q<=8'h00;
	15'h4288: q<=8'h34;
	15'h4289: q<=8'h32;
	15'h428a: q<=8'h3e;
	15'h428b: q<=8'h38;
	15'h428c: q<=8'h00;
	15'h428d: q<=8'h1a;
	15'h428e: q<=8'h24;
	15'h428f: q<=8'h16;
	15'h4290: q<=8'h30;
	15'h4291: q<=8'h22;
	15'h4292: q<=8'h1e;
	15'h4293: q<=8'hb8;
	15'h4294: q<=8'hb5;
	15'h4295: q<=8'h2a;
	15'h4296: q<=8'h30;
	15'h4297: q<=8'h32;
	15'h4298: q<=8'h34;
	15'h4299: q<=8'h20;
	15'h429a: q<=8'h00;
	15'h429b: q<=8'h1c;
	15'h429c: q<=8'h38;
	15'h429d: q<=8'h1e;
	15'h429e: q<=8'h24;
	15'h429f: q<=8'h1e;
	15'h42a0: q<=8'h30;
	15'h42a1: q<=8'h00;
	15'h42a2: q<=8'h48;
	15'h42a3: q<=8'h3e;
	15'h42a4: q<=8'h2e;
	15'h42a5: q<=8'h00;
	15'h42a6: q<=8'h42;
	15'h42a7: q<=8'h1e;
	15'h42a8: q<=8'h1a;
	15'h42a9: q<=8'h24;
	15'h42aa: q<=8'h3a;
	15'h42ab: q<=8'h1e;
	15'h42ac: q<=8'h2c;
	15'h42ad: q<=8'hb0;
	15'h42ae: q<=8'hac;
	15'h42af: q<=8'h22;
	15'h42b0: q<=8'h26;
	15'h42b1: q<=8'h38;
	15'h42b2: q<=8'h1e;
	15'h42b3: q<=8'h00;
	15'h42b4: q<=8'h2c;
	15'h42b5: q<=8'h16;
	15'h42b6: q<=8'h00;
	15'h42b7: q<=8'h34;
	15'h42b8: q<=8'h1e;
	15'h42b9: q<=8'h38;
	15'h42ba: q<=8'h26;
	15'h42bb: q<=8'h2c;
	15'h42bc: q<=8'h2c;
	15'h42bd: q<=8'h16;
	15'h42be: q<=8'h00;
	15'h42bf: q<=8'h34;
	15'h42c0: q<=8'h16;
	15'h42c1: q<=8'h38;
	15'h42c2: q<=8'h16;
	15'h42c3: q<=8'h00;
	15'h42c4: q<=8'h1a;
	15'h42c5: q<=8'h16;
	15'h42c6: q<=8'h2e;
	15'h42c7: q<=8'h18;
	15'h42c8: q<=8'h26;
	15'h42c9: q<=8'h16;
	15'h42ca: q<=8'hb8;
	15'h42cb: q<=8'hc4;
	15'h42cc: q<=8'h34;
	15'h42cd: q<=8'h38;
	15'h42ce: q<=8'h1e;
	15'h42cf: q<=8'h3a;
	15'h42d0: q<=8'h3a;
	15'h42d1: q<=8'h00;
	15'h42d2: q<=8'h20;
	15'h42d3: q<=8'h26;
	15'h42d4: q<=8'h38;
	15'h42d5: q<=8'h1e;
	15'h42d6: q<=8'h00;
	15'h42d7: q<=8'h3c;
	15'h42d8: q<=8'h32;
	15'h42d9: q<=8'h00;
	15'h42da: q<=8'h3a;
	15'h42db: q<=8'h1e;
	15'h42dc: q<=8'h2c;
	15'h42dd: q<=8'h1e;
	15'h42de: q<=8'h1a;
	15'h42df: q<=8'hbc;
	15'h42e0: q<=8'hb2;
	15'h42e1: q<=8'h34;
	15'h42e2: q<=8'h32;
	15'h42e3: q<=8'h3e;
	15'h42e4: q<=8'h3a;
	15'h42e5: q<=8'h3a;
	15'h42e6: q<=8'h1e;
	15'h42e7: q<=8'h48;
	15'h42e8: q<=8'h00;
	15'h42e9: q<=8'h20;
	15'h42ea: q<=8'h1e;
	15'h42eb: q<=8'h3e;
	15'h42ec: q<=8'h00;
	15'h42ed: q<=8'h36;
	15'h42ee: q<=8'h3e;
	15'h42ef: q<=8'h16;
	15'h42f0: q<=8'h30;
	15'h42f1: q<=8'h1c;
	15'h42f2: q<=8'h00;
	15'h42f3: q<=8'h1a;
	15'h42f4: q<=8'h32;
	15'h42f5: q<=8'h38;
	15'h42f6: q<=8'h38;
	15'h42f7: q<=8'h1e;
	15'h42f8: q<=8'h1a;
	15'h42f9: q<=8'h3c;
	15'h42fa: q<=8'h9e;
	15'h42fb: q<=8'hb2;
	15'h42fc: q<=8'h20;
	15'h42fd: q<=8'h26;
	15'h42fe: q<=8'h38;
	15'h42ff: q<=8'h1e;
	15'h4300: q<=8'h00;
	15'h4301: q<=8'h1c;
	15'h4302: q<=8'h38;
	15'h4303: q<=8'h3e;
	15'h4304: q<=8'h1e;
	15'h4305: q<=8'h1a;
	15'h4306: q<=8'h2a;
	15'h4307: q<=8'h1e;
	15'h4308: q<=8'h30;
	15'h4309: q<=8'h00;
	15'h430a: q<=8'h42;
	15'h430b: q<=8'h1e;
	15'h430c: q<=8'h30;
	15'h430d: q<=8'h30;
	15'h430e: q<=8'h00;
	15'h430f: q<=8'h38;
	15'h4310: q<=8'h26;
	15'h4311: q<=8'h1a;
	15'h4312: q<=8'h24;
	15'h4313: q<=8'h3c;
	15'h4314: q<=8'h26;
	15'h4315: q<=8'ha2;
	15'h4316: q<=8'hac;
	15'h4317: q<=8'h32;
	15'h4318: q<=8'h34;
	15'h4319: q<=8'h38;
	15'h431a: q<=8'h26;
	15'h431b: q<=8'h2e;
	15'h431c: q<=8'h16;
	15'h431d: q<=8'h00;
	15'h431e: q<=8'h20;
	15'h431f: q<=8'h26;
	15'h4320: q<=8'h38;
	15'h4321: q<=8'h1e;
	15'h4322: q<=8'h00;
	15'h4323: q<=8'h34;
	15'h4324: q<=8'h16;
	15'h4325: q<=8'h38;
	15'h4326: q<=8'h16;
	15'h4327: q<=8'h00;
	15'h4328: q<=8'h3a;
	15'h4329: q<=8'h1e;
	15'h432a: q<=8'h2c;
	15'h432b: q<=8'h1e;
	15'h432c: q<=8'h1a;
	15'h432d: q<=8'h1a;
	15'h432e: q<=8'h26;
	15'h432f: q<=8'h32;
	15'h4330: q<=8'h30;
	15'h4331: q<=8'h16;
	15'h4332: q<=8'hb8;
	15'h4333: q<=8'hbc;
	15'h4334: q<=8'h24;
	15'h4335: q<=8'h26;
	15'h4336: q<=8'h22;
	15'h4337: q<=8'h24;
	15'h4338: q<=8'h00;
	15'h4339: q<=8'h3a;
	15'h433a: q<=8'h1a;
	15'h433b: q<=8'h32;
	15'h433c: q<=8'h38;
	15'h433d: q<=8'h1e;
	15'h433e: q<=8'hba;
	15'h433f: q<=8'h9e;
	15'h4340: q<=8'h2e;
	15'h4341: q<=8'h1e;
	15'h4342: q<=8'h26;
	15'h4343: q<=8'h2c;
	15'h4344: q<=8'h2c;
	15'h4345: q<=8'h1e;
	15'h4346: q<=8'h3e;
	15'h4347: q<=8'h38;
	15'h4348: q<=8'h3a;
	15'h4349: q<=8'h00;
	15'h434a: q<=8'h3a;
	15'h434b: q<=8'h1a;
	15'h434c: q<=8'h32;
	15'h434d: q<=8'h38;
	15'h434e: q<=8'h1e;
	15'h434f: q<=8'hba;
	15'h4350: q<=8'hb0;
	15'h4351: q<=8'h24;
	15'h4352: q<=8'h32;
	15'h4353: q<=8'h1e;
	15'h4354: q<=8'h1a;
	15'h4355: q<=8'h24;
	15'h4356: q<=8'h3a;
	15'h4357: q<=8'h3c;
	15'h4358: q<=8'h48;
	15'h4359: q<=8'h16;
	15'h435a: q<=8'h24;
	15'h435b: q<=8'h2c;
	15'h435c: q<=8'h1e;
	15'h435d: q<=8'hb0;
	15'h435e: q<=8'hd4;
	15'h435f: q<=8'h38;
	15'h4360: q<=8'h1e;
	15'h4361: q<=8'h1a;
	15'h4362: q<=8'h32;
	15'h4363: q<=8'h38;
	15'h4364: q<=8'h1c;
	15'h4365: q<=8'hba;
	15'h4366: q<=8'hc2;
	15'h4367: q<=8'h38;
	15'h4368: q<=8'h16;
	15'h4369: q<=8'h30;
	15'h436a: q<=8'h2a;
	15'h436b: q<=8'h26;
	15'h436c: q<=8'h30;
	15'h436d: q<=8'h22;
	15'h436e: q<=8'h00;
	15'h436f: q<=8'h20;
	15'h4370: q<=8'h38;
	15'h4371: q<=8'h32;
	15'h4372: q<=8'h2e;
	15'h4373: q<=8'h00;
	15'h4374: q<=8'h04;
	15'h4375: q<=8'h00;
	15'h4376: q<=8'h3c;
	15'h4377: q<=8'h32;
	15'h4378: q<=8'h80;
	15'h4379: q<=8'hc2;
	15'h437a: q<=8'h34;
	15'h437b: q<=8'h2c;
	15'h437c: q<=8'h16;
	15'h437d: q<=8'h1a;
	15'h437e: q<=8'h1e;
	15'h437f: q<=8'h2e;
	15'h4380: q<=8'h1e;
	15'h4381: q<=8'h30;
	15'h4382: q<=8'h3c;
	15'h4383: q<=8'h00;
	15'h4384: q<=8'h1c;
	15'h4385: q<=8'h1e;
	15'h4386: q<=8'h00;
	15'h4387: q<=8'h04;
	15'h4388: q<=8'h00;
	15'h4389: q<=8'h16;
	15'h438a: q<=8'h80;
	15'h438b: q<=8'hbc;
	15'h438c: q<=8'h38;
	15'h438d: q<=8'h16;
	15'h438e: q<=8'h30;
	15'h438f: q<=8'h22;
	15'h4390: q<=8'h2c;
	15'h4391: q<=8'h26;
	15'h4392: q<=8'h3a;
	15'h4393: q<=8'h3c;
	15'h4394: q<=8'h1e;
	15'h4395: q<=8'h00;
	15'h4396: q<=8'h40;
	15'h4397: q<=8'h32;
	15'h4398: q<=8'h30;
	15'h4399: q<=8'h00;
	15'h439a: q<=8'h04;
	15'h439b: q<=8'h00;
	15'h439c: q<=8'h48;
	15'h439d: q<=8'h3e;
	15'h439e: q<=8'h2e;
	15'h439f: q<=8'h80;
	15'h43a0: q<=8'hc8;
	15'h43a1: q<=8'h38;
	15'h43a2: q<=8'h16;
	15'h43a3: q<=8'h30;
	15'h43a4: q<=8'h2a;
	15'h43a5: q<=8'h26;
	15'h43a6: q<=8'h30;
	15'h43a7: q<=8'h22;
	15'h43a8: q<=8'h00;
	15'h43a9: q<=8'h1c;
	15'h43aa: q<=8'h1e;
	15'h43ab: q<=8'h00;
	15'h43ac: q<=8'h04;
	15'h43ad: q<=8'h00;
	15'h43ae: q<=8'h16;
	15'h43af: q<=8'h80;
	15'h43b0: q<=8'hd9;
	15'h43b1: q<=8'h38;
	15'h43b2: q<=8'h16;
	15'h43b3: q<=8'h3c;
	15'h43b4: q<=8'h1e;
	15'h43b5: q<=8'h00;
	15'h43b6: q<=8'h46;
	15'h43b7: q<=8'h32;
	15'h43b8: q<=8'h3e;
	15'h43b9: q<=8'h38;
	15'h43ba: q<=8'h3a;
	15'h43bb: q<=8'h1e;
	15'h43bc: q<=8'h2c;
	15'h43bd: q<=8'ha0;
	15'h43be: q<=8'hdc;
	15'h43bf: q<=8'h1e;
	15'h43c0: q<=8'h40;
	15'h43c1: q<=8'h16;
	15'h43c2: q<=8'h2c;
	15'h43c3: q<=8'h3e;
	15'h43c4: q<=8'h1e;
	15'h43c5: q<=8'h48;
	15'h43c6: q<=8'h4c;
	15'h43c7: q<=8'h40;
	15'h43c8: q<=8'h32;
	15'h43c9: q<=8'h3e;
	15'h43ca: q<=8'hba;
	15'h43cb: q<=8'hd6;
	15'h43cc: q<=8'h3a;
	15'h43cd: q<=8'h1e;
	15'h43ce: q<=8'h2c;
	15'h43cf: q<=8'h18;
	15'h43d0: q<=8'h3a;
	15'h43d1: q<=8'h3c;
	15'h43d2: q<=8'h00;
	15'h43d3: q<=8'h38;
	15'h43d4: q<=8'h1e;
	15'h43d5: q<=8'h1a;
	15'h43d6: q<=8'h24;
	15'h43d7: q<=8'h30;
	15'h43d8: q<=8'h1e;
	15'h43d9: q<=8'hb0;
	15'h43da: q<=8'hdf;
	15'h43db: q<=8'h1a;
	15'h43dc: q<=8'h16;
	15'h43dd: q<=8'h2c;
	15'h43de: q<=8'h26;
	15'h43df: q<=8'h20;
	15'h43e0: q<=8'h26;
	15'h43e1: q<=8'h36;
	15'h43e2: q<=8'h3e;
	15'h43e3: q<=8'h1e;
	15'h43e4: q<=8'h3a;
	15'h43e5: q<=8'h9e;
	15'h43e6: q<=8'haa;
	15'h43e7: q<=8'h30;
	15'h43e8: q<=8'h32;
	15'h43e9: q<=8'h40;
	15'h43ea: q<=8'h26;
	15'h43eb: q<=8'h1a;
	15'h43ec: q<=8'h9e;
	15'h43ed: q<=8'haa;
	15'h43ee: q<=8'h30;
	15'h43ef: q<=8'h32;
	15'h43f0: q<=8'h40;
	15'h43f1: q<=8'h26;
	15'h43f2: q<=8'h1a;
	15'h43f3: q<=8'h26;
	15'h43f4: q<=8'hb2;
	15'h43f5: q<=8'haa;
	15'h43f6: q<=8'h16;
	15'h43f7: q<=8'h30;
	15'h43f8: q<=8'h20;
	15'h43f9: q<=8'h16;
	15'h43fa: q<=8'h1e;
	15'h43fb: q<=8'h30;
	15'h43fc: q<=8'h22;
	15'h43fd: q<=8'h1e;
	15'h43fe: q<=8'hb8;
	15'h43ff: q<=8'h4a;
	15'h4400: q<=8'h1e;
	15'h4401: q<=8'h44;
	15'h4402: q<=8'h34;
	15'h4403: q<=8'h1e;
	15'h4404: q<=8'h38;
	15'h4405: q<=8'hbc;
	15'h4406: q<=8'h45;
	15'h4407: q<=8'h1e;
	15'h4408: q<=8'h44;
	15'h4409: q<=8'h34;
	15'h440a: q<=8'h1e;
	15'h440b: q<=8'h38;
	15'h440c: q<=8'h3c;
	15'h440d: q<=8'hb2;
	15'h440e: q<=8'h40;
	15'h440f: q<=8'h1e;
	15'h4410: q<=8'h38;
	15'h4411: q<=8'h20;
	15'h4412: q<=8'h16;
	15'h4413: q<=8'h24;
	15'h4414: q<=8'h38;
	15'h4415: q<=8'h1e;
	15'h4416: q<=8'hb0;
	15'h4417: q<=8'h8b;
	15'h4418: q<=8'h18;
	15'h4419: q<=8'h32;
	15'h441a: q<=8'h30;
	15'h441b: q<=8'h3e;
	15'h441c: q<=8'hba;
	15'h441d: q<=8'he8;
	15'h441e: q<=8'h3c;
	15'h441f: q<=8'h26;
	15'h4420: q<=8'h2e;
	15'h4421: q<=8'h9e;
	15'h4422: q<=8'he0;
	15'h4423: q<=8'h1c;
	15'h4424: q<=8'h3e;
	15'h4425: q<=8'h38;
	15'h4426: q<=8'h1e;
	15'h4427: q<=8'h9e;
	15'h4428: q<=8'he8;
	15'h4429: q<=8'h48;
	15'h442a: q<=8'h1e;
	15'h442b: q<=8'h26;
	15'h442c: q<=8'hbc;
	15'h442d: q<=8'he4;
	15'h442e: q<=8'h3c;
	15'h442f: q<=8'h26;
	15'h4430: q<=8'h1e;
	15'h4431: q<=8'h2e;
	15'h4432: q<=8'h34;
	15'h4433: q<=8'hb2;
	15'h4434: q<=8'h8b;
	15'h4435: q<=8'h2c;
	15'h4436: q<=8'h1e;
	15'h4437: q<=8'h40;
	15'h4438: q<=8'h1e;
	15'h4439: q<=8'hac;
	15'h443a: q<=8'h8b;
	15'h443b: q<=8'h30;
	15'h443c: q<=8'h26;
	15'h443d: q<=8'h40;
	15'h443e: q<=8'h1e;
	15'h443f: q<=8'h16;
	15'h4440: q<=8'hbe;
	15'h4441: q<=8'h8b;
	15'h4442: q<=8'h22;
	15'h4443: q<=8'h38;
	15'h4444: q<=8'h16;
	15'h4445: q<=8'h9c;
	15'h4446: q<=8'h8b;
	15'h4447: q<=8'h30;
	15'h4448: q<=8'h26;
	15'h4449: q<=8'h40;
	15'h444a: q<=8'h1e;
	15'h444b: q<=8'hac;
	15'h444c: q<=8'h8b;
	15'h444d: q<=8'h24;
	15'h444e: q<=8'h32;
	15'h444f: q<=8'h2c;
	15'h4450: q<=8'h9e;
	15'h4451: q<=8'h8b;
	15'h4452: q<=8'h3c;
	15'h4453: q<=8'h38;
	15'h4454: q<=8'h32;
	15'h4455: q<=8'hbe;
	15'h4456: q<=8'h8b;
	15'h4457: q<=8'h24;
	15'h4458: q<=8'h32;
	15'h4459: q<=8'h46;
	15'h445a: q<=8'hb2;
	15'h445b: q<=8'h8b;
	15'h445c: q<=8'h2c;
	15'h445d: q<=8'h32;
	15'h445e: q<=8'h1a;
	15'h445f: q<=8'ha4;
	15'h4460: q<=8'hdc;
	15'h4461: q<=8'h26;
	15'h4462: q<=8'h30;
	15'h4463: q<=8'h3a;
	15'h4464: q<=8'h1e;
	15'h4465: q<=8'h38;
	15'h4466: q<=8'h3c;
	15'h4467: q<=8'h00;
	15'h4468: q<=8'h1a;
	15'h4469: q<=8'h32;
	15'h446a: q<=8'h26;
	15'h446b: q<=8'h30;
	15'h446c: q<=8'hba;
	15'h446d: q<=8'hc1;
	15'h446e: q<=8'h26;
	15'h446f: q<=8'h30;
	15'h4470: q<=8'h3c;
	15'h4471: q<=8'h38;
	15'h4472: q<=8'h32;
	15'h4473: q<=8'h1c;
	15'h4474: q<=8'h3e;
	15'h4475: q<=8'h26;
	15'h4476: q<=8'h38;
	15'h4477: q<=8'h1e;
	15'h4478: q<=8'h00;
	15'h4479: q<=8'h2c;
	15'h447a: q<=8'h1e;
	15'h447b: q<=8'h3a;
	15'h447c: q<=8'h00;
	15'h447d: q<=8'h34;
	15'h447e: q<=8'h26;
	15'h447f: q<=8'h1e;
	15'h4480: q<=8'h1a;
	15'h4481: q<=8'h1e;
	15'h4482: q<=8'hba;
	15'h4483: q<=8'hd6;
	15'h4484: q<=8'h22;
	15'h4485: q<=8'h1e;
	15'h4486: q<=8'h2c;
	15'h4487: q<=8'h1c;
	15'h4488: q<=8'h00;
	15'h4489: q<=8'h1e;
	15'h448a: q<=8'h26;
	15'h448b: q<=8'h30;
	15'h448c: q<=8'h42;
	15'h448d: q<=8'h1e;
	15'h448e: q<=8'h38;
	15'h448f: q<=8'h20;
	15'h4490: q<=8'h1e;
	15'h4491: q<=8'hb0;
	15'h4492: q<=8'hd6;
	15'h4493: q<=8'h26;
	15'h4494: q<=8'h30;
	15'h4495: q<=8'h3a;
	15'h4496: q<=8'h1e;
	15'h4497: q<=8'h38;
	15'h4498: q<=8'h3c;
	15'h4499: q<=8'h1e;
	15'h449a: q<=8'h00;
	15'h449b: q<=8'h20;
	15'h449c: q<=8'h26;
	15'h449d: q<=8'h1a;
	15'h449e: q<=8'h24;
	15'h449f: q<=8'h16;
	15'h44a0: q<=8'hba;
	15'h44a1: q<=8'h00;
	15'h44a2: q<=8'h20;
	15'h44a3: q<=8'h38;
	15'h44a4: q<=8'h1e;
	15'h44a5: q<=8'h1e;
	15'h44a6: q<=8'h00;
	15'h44a7: q<=8'h34;
	15'h44a8: q<=8'h2c;
	15'h44a9: q<=8'h16;
	15'h44aa: q<=8'hc6;
	15'h44ab: q<=8'h0e;
	15'h44ac: q<=8'h04;
	15'h44ad: q<=8'h00;
	15'h44ae: q<=8'h1a;
	15'h44af: q<=8'h32;
	15'h44b0: q<=8'h26;
	15'h44b1: q<=8'h30;
	15'h44b2: q<=8'h00;
	15'h44b3: q<=8'h06;
	15'h44b4: q<=8'h00;
	15'h44b5: q<=8'h34;
	15'h44b6: q<=8'h2c;
	15'h44b7: q<=8'h16;
	15'h44b8: q<=8'h46;
	15'h44b9: q<=8'hba;
	15'h44ba: q<=8'hfa;
	15'h44bb: q<=8'h04;
	15'h44bc: q<=8'h00;
	15'h44bd: q<=8'h34;
	15'h44be: q<=8'h26;
	15'h44bf: q<=8'h1e;
	15'h44c0: q<=8'h1a;
	15'h44c1: q<=8'h1e;
	15'h44c2: q<=8'h00;
	15'h44c3: q<=8'h06;
	15'h44c4: q<=8'h00;
	15'h44c5: q<=8'h28;
	15'h44c6: q<=8'h32;
	15'h44c7: q<=8'h3e;
	15'h44c8: q<=8'h1e;
	15'h44c9: q<=8'h3e;
	15'h44ca: q<=8'h38;
	15'h44cb: q<=8'hba;
	15'h44cc: q<=8'h00;
	15'h44cd: q<=8'h04;
	15'h44ce: q<=8'h00;
	15'h44cf: q<=8'h2e;
	15'h44d0: q<=8'h3e;
	15'h44d1: q<=8'h1e;
	15'h44d2: q<=8'h30;
	15'h44d3: q<=8'h48;
	15'h44d4: q<=8'h00;
	15'h44d5: q<=8'h06;
	15'h44d6: q<=8'h00;
	15'h44d7: q<=8'h3a;
	15'h44d8: q<=8'h34;
	15'h44d9: q<=8'h26;
	15'h44da: q<=8'h1e;
	15'h44db: q<=8'h2c;
	15'h44dc: q<=8'h9e;
	15'h44dd: q<=8'hfa;
	15'h44de: q<=8'h04;
	15'h44df: q<=8'h00;
	15'h44e0: q<=8'h2e;
	15'h44e1: q<=8'h32;
	15'h44e2: q<=8'h30;
	15'h44e3: q<=8'h1e;
	15'h44e4: q<=8'h1c;
	15'h44e5: q<=8'h16;
	15'h44e6: q<=8'h00;
	15'h44e7: q<=8'h06;
	15'h44e8: q<=8'h00;
	15'h44e9: q<=8'h28;
	15'h44ea: q<=8'h3e;
	15'h44eb: q<=8'h1e;
	15'h44ec: q<=8'h22;
	15'h44ed: q<=8'h32;
	15'h44ee: q<=8'hba;
	15'h44ef: q<=8'h14;
	15'h44f0: q<=8'h04;
	15'h44f1: q<=8'h00;
	15'h44f2: q<=8'h1a;
	15'h44f3: q<=8'h32;
	15'h44f4: q<=8'h26;
	15'h44f5: q<=8'h30;
	15'h44f6: q<=8'h00;
	15'h44f7: q<=8'h04;
	15'h44f8: q<=8'h00;
	15'h44f9: q<=8'h34;
	15'h44fa: q<=8'h2c;
	15'h44fb: q<=8'h16;
	15'h44fc: q<=8'hc6;
	15'h44fd: q<=8'h00;
	15'h44fe: q<=8'h04;
	15'h44ff: q<=8'h00;
	15'h4500: q<=8'h34;
	15'h4501: q<=8'h26;
	15'h4502: q<=8'h1e;
	15'h4503: q<=8'h1a;
	15'h4504: q<=8'h1e;
	15'h4505: q<=8'h00;
	15'h4506: q<=8'h04;
	15'h4507: q<=8'h00;
	15'h4508: q<=8'h28;
	15'h4509: q<=8'h32;
	15'h450a: q<=8'h3e;
	15'h450b: q<=8'h1e;
	15'h450c: q<=8'h3e;
	15'h450d: q<=8'hb8;
	15'h450e: q<=8'h00;
	15'h450f: q<=8'h04;
	15'h4510: q<=8'h00;
	15'h4511: q<=8'h2e;
	15'h4512: q<=8'h3e;
	15'h4513: q<=8'h1e;
	15'h4514: q<=8'h30;
	15'h4515: q<=8'h48;
	15'h4516: q<=8'h1e;
	15'h4517: q<=8'h00;
	15'h4518: q<=8'h04;
	15'h4519: q<=8'h00;
	15'h451a: q<=8'h3a;
	15'h451b: q<=8'h34;
	15'h451c: q<=8'h26;
	15'h451d: q<=8'h1e;
	15'h451e: q<=8'hac;
	15'h451f: q<=8'h00;
	15'h4520: q<=8'h04;
	15'h4521: q<=8'h00;
	15'h4522: q<=8'h2e;
	15'h4523: q<=8'h32;
	15'h4524: q<=8'h30;
	15'h4525: q<=8'h1e;
	15'h4526: q<=8'h1c;
	15'h4527: q<=8'h16;
	15'h4528: q<=8'h00;
	15'h4529: q<=8'h04;
	15'h452a: q<=8'h00;
	15'h452b: q<=8'h28;
	15'h452c: q<=8'h3e;
	15'h452d: q<=8'h1e;
	15'h452e: q<=8'h22;
	15'h452f: q<=8'hb2;
	15'h4530: q<=8'h0e;
	15'h4531: q<=8'h06;
	15'h4532: q<=8'h00;
	15'h4533: q<=8'h1a;
	15'h4534: q<=8'h32;
	15'h4535: q<=8'h26;
	15'h4536: q<=8'h30;
	15'h4537: q<=8'h3a;
	15'h4538: q<=8'h00;
	15'h4539: q<=8'h04;
	15'h453a: q<=8'h00;
	15'h453b: q<=8'h34;
	15'h453c: q<=8'h2c;
	15'h453d: q<=8'h16;
	15'h453e: q<=8'hc6;
	15'h453f: q<=8'hfa;
	15'h4540: q<=8'h06;
	15'h4541: q<=8'h00;
	15'h4542: q<=8'h34;
	15'h4543: q<=8'h26;
	15'h4544: q<=8'h1e;
	15'h4545: q<=8'h1a;
	15'h4546: q<=8'h1e;
	15'h4547: q<=8'h3a;
	15'h4548: q<=8'h00;
	15'h4549: q<=8'h04;
	15'h454a: q<=8'h00;
	15'h454b: q<=8'h28;
	15'h454c: q<=8'h32;
	15'h454d: q<=8'h3e;
	15'h454e: q<=8'h1e;
	15'h454f: q<=8'h3e;
	15'h4550: q<=8'hb8;
	15'h4551: q<=8'hfa;
	15'h4552: q<=8'h06;
	15'h4553: q<=8'h00;
	15'h4554: q<=8'h2e;
	15'h4555: q<=8'h3e;
	15'h4556: q<=8'h1e;
	15'h4557: q<=8'h30;
	15'h4558: q<=8'h48;
	15'h4559: q<=8'h1e;
	15'h455a: q<=8'h30;
	15'h455b: q<=8'h00;
	15'h455c: q<=8'h04;
	15'h455d: q<=8'h00;
	15'h455e: q<=8'h3a;
	15'h455f: q<=8'h34;
	15'h4560: q<=8'h26;
	15'h4561: q<=8'h1e;
	15'h4562: q<=8'hac;
	15'h4563: q<=8'hfa;
	15'h4564: q<=8'h06;
	15'h4565: q<=8'h00;
	15'h4566: q<=8'h2e;
	15'h4567: q<=8'h32;
	15'h4568: q<=8'h30;
	15'h4569: q<=8'h1e;
	15'h456a: q<=8'h1c;
	15'h456b: q<=8'h16;
	15'h456c: q<=8'h3a;
	15'h456d: q<=8'h00;
	15'h456e: q<=8'h04;
	15'h456f: q<=8'h00;
	15'h4570: q<=8'h28;
	15'h4571: q<=8'h3e;
	15'h4572: q<=8'h1e;
	15'h4573: q<=8'h22;
	15'h4574: q<=8'hb2;
	15'h4575: q<=8'hd3;
	15'h4576: q<=8'h50;
	15'h4577: q<=8'h00;
	15'h4578: q<=8'h2e;
	15'h4579: q<=8'h1a;
	15'h457a: q<=8'h2e;
	15'h457b: q<=8'h2c;
	15'h457c: q<=8'h44;
	15'h457d: q<=8'h44;
	15'h457e: q<=8'h44;
	15'h457f: q<=8'h00;
	15'h4580: q<=8'h16;
	15'h4581: q<=8'h3c;
	15'h4582: q<=8'h16;
	15'h4583: q<=8'h38;
	15'h4584: q<=8'ha6;
	15'h4585: q<=8'ha0;
	15'h4586: q<=8'h1a;
	15'h4587: q<=8'h38;
	15'h4588: q<=8'h1e;
	15'h4589: q<=8'h1c;
	15'h458a: q<=8'h26;
	15'h458b: q<=8'h3c;
	15'h458c: q<=8'h3a;
	15'h458d: q<=8'h80;
	15'h458e: q<=8'ha0;
	15'h458f: q<=8'h2a;
	15'h4590: q<=8'h38;
	15'h4591: q<=8'h1e;
	15'h4592: q<=8'h1c;
	15'h4593: q<=8'h26;
	15'h4594: q<=8'h3c;
	15'h4595: q<=8'h1e;
	15'h4596: q<=8'h80;
	15'h4597: q<=8'ha0;
	15'h4598: q<=8'h1a;
	15'h4599: q<=8'h38;
	15'h459a: q<=8'h1e;
	15'h459b: q<=8'h1c;
	15'h459c: q<=8'h26;
	15'h459d: q<=8'h3c;
	15'h459e: q<=8'h32;
	15'h459f: q<=8'h3a;
	15'h45a0: q<=8'h80;
	15'h45a1: q<=8'hda;
	15'h45a2: q<=8'h18;
	15'h45a3: q<=8'h32;
	15'h45a4: q<=8'h30;
	15'h45a5: q<=8'h3e;
	15'h45a6: q<=8'h3a;
	15'h45a7: q<=8'h80;
	15'h45a8: q<=8'hd0;
	15'h45a9: q<=8'h06;
	15'h45aa: q<=8'h00;
	15'h45ab: q<=8'h1a;
	15'h45ac: q<=8'h38;
	15'h45ad: q<=8'h1e;
	15'h45ae: q<=8'h1c;
	15'h45af: q<=8'h26;
	15'h45b0: q<=8'h3c;
	15'h45b1: q<=8'h00;
	15'h45b2: q<=8'h2e;
	15'h45b3: q<=8'h26;
	15'h45b4: q<=8'h30;
	15'h45b5: q<=8'h26;
	15'h45b6: q<=8'h2e;
	15'h45b7: q<=8'h3e;
	15'h45b8: q<=8'hae;
	15'h45b9: q<=8'hd6;
	15'h45ba: q<=8'h06;
	15'h45bb: q<=8'h00;
	15'h45bc: q<=8'h28;
	15'h45bd: q<=8'h1e;
	15'h45be: q<=8'h3e;
	15'h45bf: q<=8'h44;
	15'h45c0: q<=8'h00;
	15'h45c1: q<=8'h2e;
	15'h45c2: q<=8'h26;
	15'h45c3: q<=8'h30;
	15'h45c4: q<=8'h26;
	15'h45c5: q<=8'h2e;
	15'h45c6: q<=8'h3e;
	15'h45c7: q<=8'hae;
	15'h45c8: q<=8'hd0;
	15'h45c9: q<=8'h06;
	15'h45ca: q<=8'h00;
	15'h45cb: q<=8'h3a;
	15'h45cc: q<=8'h34;
	15'h45cd: q<=8'h26;
	15'h45ce: q<=8'h1e;
	15'h45cf: q<=8'h2c;
	15'h45d0: q<=8'h1e;
	15'h45d1: q<=8'h00;
	15'h45d2: q<=8'h2e;
	15'h45d3: q<=8'h26;
	15'h45d4: q<=8'h30;
	15'h45d5: q<=8'h26;
	15'h45d6: q<=8'h2e;
	15'h45d7: q<=8'h3e;
	15'h45d8: q<=8'hae;
	15'h45d9: q<=8'hd3;
	15'h45da: q<=8'h06;
	15'h45db: q<=8'h00;
	15'h45dc: q<=8'h28;
	15'h45dd: q<=8'h3e;
	15'h45de: q<=8'h1e;
	15'h45df: q<=8'h22;
	15'h45e0: q<=8'h32;
	15'h45e1: q<=8'h3a;
	15'h45e2: q<=8'h00;
	15'h45e3: q<=8'h2e;
	15'h45e4: q<=8'h26;
	15'h45e5: q<=8'h30;
	15'h45e6: q<=8'h26;
	15'h45e7: q<=8'h2e;
	15'h45e8: q<=8'hb2;
	15'h45e9: q<=8'hc8;
	15'h45ea: q<=8'h18;
	15'h45eb: q<=8'h32;
	15'h45ec: q<=8'h30;
	15'h45ed: q<=8'h3e;
	15'h45ee: q<=8'h3a;
	15'h45ef: q<=8'h00;
	15'h45f0: q<=8'h1e;
	15'h45f1: q<=8'h40;
	15'h45f2: q<=8'h1e;
	15'h45f3: q<=8'h38;
	15'h45f4: q<=8'h46;
	15'h45f5: q<=8'h80;
	15'h45f6: q<=8'hce;
	15'h45f7: q<=8'h18;
	15'h45f8: q<=8'h32;
	15'h45f9: q<=8'h30;
	15'h45fa: q<=8'h3e;
	15'h45fb: q<=8'h3a;
	15'h45fc: q<=8'h00;
	15'h45fd: q<=8'h1a;
	15'h45fe: q<=8'h24;
	15'h45ff: q<=8'h16;
	15'h4600: q<=8'h36;
	15'h4601: q<=8'h3e;
	15'h4602: q<=8'h1e;
	15'h4603: q<=8'h80;
	15'h4604: q<=8'hce;
	15'h4605: q<=8'h18;
	15'h4606: q<=8'h32;
	15'h4607: q<=8'h30;
	15'h4608: q<=8'h3e;
	15'h4609: q<=8'h3a;
	15'h460a: q<=8'h00;
	15'h460b: q<=8'h28;
	15'h460c: q<=8'h1e;
	15'h460d: q<=8'h1c;
	15'h460e: q<=8'h1e;
	15'h460f: q<=8'h80;
	15'h4610: q<=8'hc8;
	15'h4611: q<=8'h18;
	15'h4612: q<=8'h32;
	15'h4613: q<=8'h30;
	15'h4614: q<=8'h3e;
	15'h4615: q<=8'h3a;
	15'h4616: q<=8'h00;
	15'h4617: q<=8'h1a;
	15'h4618: q<=8'h16;
	15'h4619: q<=8'h1c;
	15'h461a: q<=8'h16;
	15'h461b: q<=8'h80;
	15'h461c: q<=8'hb8;
	15'h461d: q<=8'h16;
	15'h461e: q<=8'h40;
	15'h461f: q<=8'h32;
	15'h4620: q<=8'h26;
	15'h4621: q<=8'h1c;
	15'h4622: q<=8'h00;
	15'h4623: q<=8'h3a;
	15'h4624: q<=8'h34;
	15'h4625: q<=8'h26;
	15'h4626: q<=8'h2a;
	15'h4627: q<=8'h1e;
	15'h4628: q<=8'hba;
	15'h4629: q<=8'h88;
	15'h462a: q<=8'h16;
	15'h462b: q<=8'h3c;
	15'h462c: q<=8'h3c;
	15'h462d: q<=8'h1e;
	15'h462e: q<=8'h30;
	15'h462f: q<=8'h3c;
	15'h4630: q<=8'h26;
	15'h4631: q<=8'h32;
	15'h4632: q<=8'h30;
	15'h4633: q<=8'h00;
	15'h4634: q<=8'h16;
	15'h4635: q<=8'h3e;
	15'h4636: q<=8'h44;
	15'h4637: q<=8'h00;
	15'h4638: q<=8'h2c;
	15'h4639: q<=8'h16;
	15'h463a: q<=8'h30;
	15'h463b: q<=8'h1a;
	15'h463c: q<=8'h1e;
	15'h463d: q<=8'hba;
	15'h463e: q<=8'h96;
	15'h463f: q<=8'h3a;
	15'h4640: q<=8'h34;
	15'h4641: q<=8'h26;
	15'h4642: q<=8'h3c;
	15'h4643: q<=8'h48;
	15'h4644: q<=8'h1e;
	15'h4645: q<=8'h30;
	15'h4646: q<=8'h00;
	15'h4647: q<=8'h16;
	15'h4648: q<=8'h3e;
	15'h4649: q<=8'h3a;
	15'h464a: q<=8'h42;
	15'h464b: q<=8'h1e;
	15'h464c: q<=8'h26;
	15'h464d: q<=8'h1a;
	15'h464e: q<=8'h24;
	15'h464f: q<=8'h1e;
	15'h4650: q<=8'hb0;
	15'h4651: q<=8'ha0;
	15'h4652: q<=8'h1e;
	15'h4653: q<=8'h40;
	15'h4654: q<=8'h26;
	15'h4655: q<=8'h3c;
	15'h4656: q<=8'h1e;
	15'h4657: q<=8'h00;
	15'h4658: q<=8'h2c;
	15'h4659: q<=8'h16;
	15'h465a: q<=8'h3a;
	15'h465b: q<=8'h00;
	15'h465c: q<=8'h34;
	15'h465d: q<=8'h3e;
	15'h465e: q<=8'h30;
	15'h465f: q<=8'h3c;
	15'h4660: q<=8'h16;
	15'h4661: q<=8'hba;
	15'h4662: q<=8'he0;
	15'h4663: q<=8'h2c;
	15'h4664: q<=8'h1e;
	15'h4665: q<=8'h40;
	15'h4666: q<=8'h1e;
	15'h4667: q<=8'hac;
	15'h4668: q<=8'hda;
	15'h4669: q<=8'h30;
	15'h466a: q<=8'h26;
	15'h466b: q<=8'h40;
	15'h466c: q<=8'h1e;
	15'h466d: q<=8'h16;
	15'h466e: q<=8'hbe;
	15'h466f: q<=8'he2;
	15'h4670: q<=8'h22;
	15'h4671: q<=8'h38;
	15'h4672: q<=8'h16;
	15'h4673: q<=8'h9c;
	15'h4674: q<=8'he0;
	15'h4675: q<=8'h30;
	15'h4676: q<=8'h26;
	15'h4677: q<=8'h40;
	15'h4678: q<=8'h1e;
	15'h4679: q<=8'hac;
	15'h467a: q<=8'hc4;
	15'h467b: q<=8'h3a;
	15'h467c: q<=8'h3e;
	15'h467d: q<=8'h34;
	15'h467e: q<=8'h1e;
	15'h467f: q<=8'h38;
	15'h4680: q<=8'h48;
	15'h4681: q<=8'h16;
	15'h4682: q<=8'h34;
	15'h4683: q<=8'h34;
	15'h4684: q<=8'h1e;
	15'h4685: q<=8'h38;
	15'h4686: q<=8'h00;
	15'h4687: q<=8'h38;
	15'h4688: q<=8'h1e;
	15'h4689: q<=8'h1a;
	15'h468a: q<=8'h24;
	15'h468b: q<=8'h16;
	15'h468c: q<=8'h38;
	15'h468d: q<=8'h22;
	15'h468e: q<=8'h9e;
	15'h468f: q<=8'hcd;
	15'h4690: q<=8'h30;
	15'h4691: q<=8'h1e;
	15'h4692: q<=8'h3e;
	15'h4693: q<=8'h1e;
	15'h4694: q<=8'h38;
	15'h4695: q<=8'h00;
	15'h4696: q<=8'h3a;
	15'h4697: q<=8'h3e;
	15'h4698: q<=8'h34;
	15'h4699: q<=8'h1e;
	15'h469a: q<=8'h38;
	15'h469b: q<=8'h48;
	15'h469c: q<=8'h16;
	15'h469d: q<=8'h34;
	15'h469e: q<=8'h34;
	15'h469f: q<=8'h1e;
	15'h46a0: q<=8'hb8;
	15'h46a1: q<=8'hcd;
	15'h46a2: q<=8'h30;
	15'h46a3: q<=8'h3e;
	15'h46a4: q<=8'h1e;
	15'h46a5: q<=8'h40;
	15'h46a6: q<=8'h32;
	15'h46a7: q<=8'h00;
	15'h46a8: q<=8'h3a;
	15'h46a9: q<=8'h3e;
	15'h46aa: q<=8'h34;
	15'h46ab: q<=8'h1e;
	15'h46ac: q<=8'h38;
	15'h46ad: q<=8'h48;
	15'h46ae: q<=8'h16;
	15'h46af: q<=8'h34;
	15'h46b0: q<=8'h34;
	15'h46b1: q<=8'h1e;
	15'h46b2: q<=8'hb8;
	15'h46b3: q<=8'h31;
	15'h46b4: q<=8'hd0;
	15'h46b5: q<=8'h6d;
	15'h46b6: q<=8'hd0;
	15'h46b7: q<=8'ha9;
	15'h46b8: q<=8'hd0;
	15'h46b9: q<=8'he5;
	15'h46ba: q<=8'hd0;
	15'h46bb: q<=8'had;
	15'h46bc: q<=8'h00;
	15'h46bd: q<=8'h0e;
	15'h46be: q<=8'h85;
	15'h46bf: q<=8'h0a;
	15'h46c0: q<=8'h29;
	15'h46c1: q<=8'h38;
	15'h46c2: q<=8'h4a;
	15'h46c3: q<=8'h4a;
	15'h46c4: q<=8'h4a;
	15'h46c5: q<=8'haa;
	15'h46c6: q<=8'hbd;
	15'h46c7: q<=8'hf7;
	15'h46c8: q<=8'hd6;
	15'h46c9: q<=8'h8d;
	15'h46ca: q<=8'h56;
	15'h46cb: q<=8'h01;
	15'h46cc: q<=8'had;
	15'h46cd: q<=8'h00;
	15'h46ce: q<=8'h0d;
	15'h46cf: q<=8'h49;
	15'h46d0: q<=8'h02;
	15'h46d1: q<=8'h85;
	15'h46d2: q<=8'h09;
	15'h46d3: q<=8'ha5;
	15'h46d4: q<=8'h0a;
	15'h46d5: q<=8'h2a;
	15'h46d6: q<=8'h2a;
	15'h46d7: q<=8'h2a;
	15'h46d8: q<=8'h29;
	15'h46d9: q<=8'h03;
	15'h46da: q<=8'haa;
	15'h46db: q<=8'hbd;
	15'h46dc: q<=8'hff;
	15'h46dd: q<=8'hd6;
	15'h46de: q<=8'h8d;
	15'h46df: q<=8'h58;
	15'h46e0: q<=8'h01;
	15'h46e1: q<=8'ha5;
	15'h46e2: q<=8'h0a;
	15'h46e3: q<=8'h29;
	15'h46e4: q<=8'h06;
	15'h46e5: q<=8'ha8;
	15'h46e6: q<=8'hb9;
	15'h46e7: q<=8'hb3;
	15'h46e8: q<=8'hd6;
	15'h46e9: q<=8'h85;
	15'h46ea: q<=8'hac;
	15'h46eb: q<=8'hb9;
	15'h46ec: q<=8'hb4;
	15'h46ed: q<=8'hd6;
	15'h46ee: q<=8'h85;
	15'h46ef: q<=8'had;
	15'h46f0: q<=8'h20;
	15'h46f1: q<=8'he0;
	15'h46f2: q<=8'hdb;
	15'h46f3: q<=8'h8d;
	15'h46f4: q<=8'h6a;
	15'h46f5: q<=8'h01;
	15'h46f6: q<=8'h60;
	15'h46f7: q<=8'h02;
	15'h46f8: q<=8'h01;
	15'h46f9: q<=8'h03;
	15'h46fa: q<=8'h04;
	15'h46fb: q<=8'h05;
	15'h46fc: q<=8'h06;
	15'h46fd: q<=8'h07;
	15'h46fe: q<=8'h00;
	15'h46ff: q<=8'h03;
	15'h4700: q<=8'h04;
	15'h4701: q<=8'h05;
	15'h4702: q<=8'h02;
	15'h4703: q<=8'h7c;
	15'h4704: q<=8'h48;
	15'h4705: q<=8'h8a;
	15'h4706: q<=8'h48;
	15'h4707: q<=8'h98;
	15'h4708: q<=8'h48;
	15'h4709: q<=8'hd8;
	15'h470a: q<=8'hba;
	15'h470b: q<=8'he0;
	15'h470c: q<=8'hd0;
	15'h470d: q<=8'h90;
	15'h470e: q<=8'h04;
	15'h470f: q<=8'ha5;
	15'h4710: q<=8'h53;
	15'h4711: q<=8'h10;
	15'h4712: q<=8'h04;
	15'h4713: q<=8'h00;
	15'h4714: q<=8'h4c;
	15'h4715: q<=8'h3f;
	15'h4716: q<=8'hd9;
	15'h4717: q<=8'h8d;
	15'h4718: q<=8'h00;
	15'h4719: q<=8'h50;
	15'h471a: q<=8'h8d;
	15'h471b: q<=8'hcb;
	15'h471c: q<=8'h60;
	15'h471d: q<=8'had;
	15'h471e: q<=8'hc8;
	15'h471f: q<=8'h60;
	15'h4720: q<=8'h49;
	15'h4721: q<=8'h0f;
	15'h4722: q<=8'ha8;
	15'h4723: q<=8'h29;
	15'h4724: q<=8'h10;
	15'h4725: q<=8'h8d;
	15'h4726: q<=8'h17;
	15'h4727: q<=8'h01;
	15'h4728: q<=8'h98;
	15'h4729: q<=8'h38;
	15'h472a: q<=8'he5;
	15'h472b: q<=8'h52;
	15'h472c: q<=8'h29;
	15'h472d: q<=8'h0f;
	15'h472e: q<=8'hc9;
	15'h472f: q<=8'h08;
	15'h4730: q<=8'h90;
	15'h4731: q<=8'h02;
	15'h4732: q<=8'h09;
	15'h4733: q<=8'hf0;
	15'h4734: q<=8'h18;
	15'h4735: q<=8'h65;
	15'h4736: q<=8'h50;
	15'h4737: q<=8'h85;
	15'h4738: q<=8'h50;
	15'h4739: q<=8'h84;
	15'h473a: q<=8'h52;
	15'h473b: q<=8'h8d;
	15'h473c: q<=8'hdb;
	15'h473d: q<=8'h60;
	15'h473e: q<=8'hac;
	15'h473f: q<=8'hd8;
	15'h4740: q<=8'h60;
	15'h4741: q<=8'had;
	15'h4742: q<=8'h00;
	15'h4743: q<=8'h0c;
	15'h4744: q<=8'h85;
	15'h4745: q<=8'h08;
	15'h4746: q<=8'ha5;
	15'h4747: q<=8'h4c;
	15'h4748: q<=8'h84;
	15'h4749: q<=8'h4c;
	15'h474a: q<=8'ha8;
	15'h474b: q<=8'h25;
	15'h474c: q<=8'h4c;
	15'h474d: q<=8'h05;
	15'h474e: q<=8'h4d;
	15'h474f: q<=8'h85;
	15'h4750: q<=8'h4d;
	15'h4751: q<=8'h98;
	15'h4752: q<=8'h05;
	15'h4753: q<=8'h4c;
	15'h4754: q<=8'h25;
	15'h4755: q<=8'h4d;
	15'h4756: q<=8'h85;
	15'h4757: q<=8'h4d;
	15'h4758: q<=8'ha8;
	15'h4759: q<=8'h45;
	15'h475a: q<=8'h4f;
	15'h475b: q<=8'h25;
	15'h475c: q<=8'h4d;
	15'h475d: q<=8'h05;
	15'h475e: q<=8'h4e;
	15'h475f: q<=8'h85;
	15'h4760: q<=8'h4e;
	15'h4761: q<=8'h84;
	15'h4762: q<=8'h4f;
	15'h4763: q<=8'ha5;
	15'h4764: q<=8'hb4;
	15'h4765: q<=8'ha4;
	15'h4766: q<=8'h13;
	15'h4767: q<=8'h10;
	15'h4768: q<=8'h02;
	15'h4769: q<=8'h09;
	15'h476a: q<=8'h04;
	15'h476b: q<=8'ha4;
	15'h476c: q<=8'h14;
	15'h476d: q<=8'h10;
	15'h476e: q<=8'h02;
	15'h476f: q<=8'h09;
	15'h4770: q<=8'h02;
	15'h4771: q<=8'ha4;
	15'h4772: q<=8'h15;
	15'h4773: q<=8'h10;
	15'h4774: q<=8'h02;
	15'h4775: q<=8'h09;
	15'h4776: q<=8'h01;
	15'h4777: q<=8'h8d;
	15'h4778: q<=8'h00;
	15'h4779: q<=8'h40;
	15'h477a: q<=8'ha6;
	15'h477b: q<=8'h3e;
	15'h477c: q<=8'he8;
	15'h477d: q<=8'ha4;
	15'h477e: q<=8'h05;
	15'h477f: q<=8'hd0;
	15'h4780: q<=8'h10;
	15'h4781: q<=8'ha2;
	15'h4782: q<=8'h00;
	15'h4783: q<=8'ha4;
	15'h4784: q<=8'h07;
	15'h4785: q<=8'hc0;
	15'h4786: q<=8'h40;
	15'h4787: q<=8'h90;
	15'h4788: q<=8'h08;
	15'h4789: q<=8'ha6;
	15'h478a: q<=8'h06;
	15'h478b: q<=8'he0;
	15'h478c: q<=8'h02;
	15'h478d: q<=8'h90;
	15'h478e: q<=8'h02;
	15'h478f: q<=8'ha2;
	15'h4790: q<=8'h03;
	15'h4791: q<=8'hbd;
	15'h4792: q<=8'hdd;
	15'h4793: q<=8'hd7;
	15'h4794: q<=8'h45;
	15'h4795: q<=8'ha1;
	15'h4796: q<=8'h29;
	15'h4797: q<=8'h03;
	15'h4798: q<=8'h45;
	15'h4799: q<=8'ha1;
	15'h479a: q<=8'h85;
	15'h479b: q<=8'ha1;
	15'h479c: q<=8'h8d;
	15'h479d: q<=8'he0;
	15'h479e: q<=8'h60;
	15'h479f: q<=8'h20;
	15'h47a0: q<=8'h24;
	15'h47a1: q<=8'hcf;
	15'h47a2: q<=8'h20;
	15'h47a3: q<=8'h0a;
	15'h47a4: q<=8'hcd;
	15'h47a5: q<=8'he6;
	15'h47a6: q<=8'h53;
	15'h47a7: q<=8'he6;
	15'h47a8: q<=8'h07;
	15'h47a9: q<=8'hd0;
	15'h47aa: q<=8'h1e;
	15'h47ab: q<=8'hee;
	15'h47ac: q<=8'h06;
	15'h47ad: q<=8'h04;
	15'h47ae: q<=8'hd0;
	15'h47af: q<=8'h08;
	15'h47b0: q<=8'hee;
	15'h47b1: q<=8'h07;
	15'h47b2: q<=8'h04;
	15'h47b3: q<=8'hd0;
	15'h47b4: q<=8'h03;
	15'h47b5: q<=8'hee;
	15'h47b6: q<=8'h08;
	15'h47b7: q<=8'h04;
	15'h47b8: q<=8'h24;
	15'h47b9: q<=8'h05;
	15'h47ba: q<=8'h50;
	15'h47bb: q<=8'h0d;
	15'h47bc: q<=8'hee;
	15'h47bd: q<=8'h09;
	15'h47be: q<=8'h04;
	15'h47bf: q<=8'hd0;
	15'h47c0: q<=8'h08;
	15'h47c1: q<=8'hee;
	15'h47c2: q<=8'h0a;
	15'h47c3: q<=8'h04;
	15'h47c4: q<=8'hd0;
	15'h47c5: q<=8'h03;
	15'h47c6: q<=8'hee;
	15'h47c7: q<=8'h0b;
	15'h47c8: q<=8'h04;
	15'h47c9: q<=8'h2c;
	15'h47ca: q<=8'h00;
	15'h47cb: q<=8'h0c;
	15'h47cc: q<=8'h50;
	15'h47cd: q<=8'h09;
	15'h47ce: q<=8'hee;
	15'h47cf: q<=8'h33;
	15'h47d0: q<=8'h01;
	15'h47d1: q<=8'h8d;
	15'h47d2: q<=8'h00;
	15'h47d3: q<=8'h58;
	15'h47d4: q<=8'h8d;
	15'h47d5: q<=8'h00;
	15'h47d6: q<=8'h48;
	15'h47d7: q<=8'h68;
	15'h47d8: q<=8'ha8;
	15'h47d9: q<=8'h68;
	15'h47da: q<=8'haa;
	15'h47db: q<=8'h68;
	15'h47dc: q<=8'h40;
	15'h47dd: q<=8'hff;
	15'h47de: q<=8'hfd;
	15'h47df: q<=8'hfe;
	15'h47e0: q<=8'hfc;
	15'h47e1: q<=8'ha9;
	15'h47e2: q<=8'h00;
	15'h47e3: q<=8'h85;
	15'h47e4: q<=8'h05;
	15'h47e5: q<=8'ha9;
	15'h47e6: q<=8'h02;
	15'h47e7: q<=8'h85;
	15'h47e8: q<=8'h01;
	15'h47e9: q<=8'had;
	15'h47ea: q<=8'hca;
	15'h47eb: q<=8'h01;
	15'h47ec: q<=8'hd0;
	15'h47ed: q<=8'h15;
	15'h47ee: q<=8'had;
	15'h47ef: q<=8'h00;
	15'h47f0: q<=8'h0c;
	15'h47f1: q<=8'h29;
	15'h47f2: q<=8'h10;
	15'h47f3: q<=8'hf0;
	15'h47f4: q<=8'h0e;
	15'h47f5: q<=8'ha9;
	15'h47f6: q<=8'h00;
	15'h47f7: q<=8'h85;
	15'h47f8: q<=8'h00;
	15'h47f9: q<=8'had;
	15'h47fa: q<=8'hc9;
	15'h47fb: q<=8'h01;
	15'h47fc: q<=8'h29;
	15'h47fd: q<=8'h03;
	15'h47fe: q<=8'hf0;
	15'h47ff: q<=8'h03;
	15'h4800: q<=8'h20;
	15'h4801: q<=8'hac;
	15'h4802: q<=8'hab;
	15'h4803: q<=8'h60;
	15'h4804: q<=8'h20;
	15'h4805: q<=8'hbb;
	15'h4806: q<=8'hd6;
	15'h4807: q<=8'h20;
	15'h4808: q<=8'ha8;
	15'h4809: q<=8'haa;
	15'h480a: q<=8'h20;
	15'h480b: q<=8'h0d;
	15'h480c: q<=8'hdd;
	15'h480d: q<=8'h20;
	15'h480e: q<=8'h41;
	15'h480f: q<=8'hdd;
	15'h4810: q<=8'had;
	15'h4811: q<=8'h58;
	15'h4812: q<=8'h01;
	15'h4813: q<=8'h85;
	15'h4814: q<=8'h37;
	15'h4815: q<=8'h20;
	15'h4816: q<=8'h53;
	15'h4817: q<=8'hdf;
	15'h4818: q<=8'ha9;
	15'h4819: q<=8'he8;
	15'h481a: q<=8'ha2;
	15'h481b: q<=8'hc0;
	15'h481c: q<=8'h20;
	15'h481d: q<=8'h75;
	15'h481e: q<=8'hdf;
	15'h481f: q<=8'ha9;
	15'h4820: q<=8'h32;
	15'h4821: q<=8'ha2;
	15'h4822: q<=8'h6c;
	15'h4823: q<=8'h20;
	15'h4824: q<=8'h39;
	15'h4825: q<=8'hdf;
	15'h4826: q<=8'hc6;
	15'h4827: q<=8'h37;
	15'h4828: q<=8'hd0;
	15'h4829: q<=8'hf5;
	15'h482a: q<=8'had;
	15'h482b: q<=8'h6a;
	15'h482c: q<=8'h01;
	15'h482d: q<=8'h29;
	15'h482e: q<=8'h03;
	15'h482f: q<=8'h0a;
	15'h4830: q<=8'ha8;
	15'h4831: q<=8'hb9;
	15'h4832: q<=8'h1f;
	15'h4833: q<=8'h3f;
	15'h4834: q<=8'hbe;
	15'h4835: q<=8'h1e;
	15'h4836: q<=8'h3f;
	15'h4837: q<=8'h20;
	15'h4838: q<=8'h39;
	15'h4839: q<=8'hdf;
	15'h483a: q<=8'had;
	15'h483b: q<=8'h00;
	15'h483c: q<=8'h02;
	15'h483d: q<=8'h20;
	15'h483e: q<=8'hce;
	15'h483f: q<=8'had;
	15'h4840: q<=8'h8d;
	15'h4841: q<=8'h00;
	15'h4842: q<=8'h02;
	15'h4843: q<=8'h29;
	15'h4844: q<=8'h06;
	15'h4845: q<=8'h48;
	15'h4846: q<=8'ha8;
	15'h4847: q<=8'hb9;
	15'h4848: q<=8'h17;
	15'h4849: q<=8'h3f;
	15'h484a: q<=8'hbe;
	15'h484b: q<=8'h16;
	15'h484c: q<=8'h3f;
	15'h484d: q<=8'h20;
	15'h484e: q<=8'h39;
	15'h484f: q<=8'hdf;
	15'h4850: q<=8'h68;
	15'h4851: q<=8'h4a;
	15'h4852: q<=8'haa;
	15'h4853: q<=8'ha5;
	15'h4854: q<=8'h4d;
	15'h4855: q<=8'h3d;
	15'h4856: q<=8'hb6;
	15'h4857: q<=8'hd8;
	15'h4858: q<=8'hdd;
	15'h4859: q<=8'hb6;
	15'h485a: q<=8'hd8;
	15'h485b: q<=8'hd0;
	15'h485c: q<=8'h1a;
	15'h485d: q<=8'hca;
	15'h485e: q<=8'hca;
	15'h485f: q<=8'h10;
	15'h4860: q<=8'h03;
	15'h4861: q<=8'h4c;
	15'h4862: q<=8'h3f;
	15'h4863: q<=8'hd9;
	15'h4864: q<=8'hd0;
	15'h4865: q<=8'h06;
	15'h4866: q<=8'h20;
	15'h4867: q<=8'he9;
	15'h4868: q<=8'hdd;
	15'h4869: q<=8'hb8;
	15'h486a: q<=8'h50;
	15'h486b: q<=8'h0b;
	15'h486c: q<=8'h20;
	15'h486d: q<=8'hed;
	15'h486e: q<=8'hdd;
	15'h486f: q<=8'had;
	15'h4870: q<=8'hc9;
	15'h4871: q<=8'h01;
	15'h4872: q<=8'h09;
	15'h4873: q<=8'h03;
	15'h4874: q<=8'h8d;
	15'h4875: q<=8'hc9;
	15'h4876: q<=8'h01;
	15'h4877: q<=8'had;
	15'h4878: q<=8'hca;
	15'h4879: q<=8'h01;
	15'h487a: q<=8'h2d;
	15'h487b: q<=8'hc6;
	15'h487c: q<=8'h01;
	15'h487d: q<=8'hf0;
	15'h487e: q<=8'h07;
	15'h487f: q<=8'ha9;
	15'h4880: q<=8'h34;
	15'h4881: q<=8'ha2;
	15'h4882: q<=8'h6e;
	15'h4883: q<=8'h20;
	15'h4884: q<=8'h39;
	15'h4885: q<=8'hdf;
	15'h4886: q<=8'h20;
	15'h4887: q<=8'h53;
	15'h4888: q<=8'hdf;
	15'h4889: q<=8'ha5;
	15'h488a: q<=8'h09;
	15'h488b: q<=8'h29;
	15'h488c: q<=8'h1c;
	15'h488d: q<=8'h4a;
	15'h488e: q<=8'h4a;
	15'h488f: q<=8'haa;
	15'h4890: q<=8'hbd;
	15'h4891: q<=8'hba;
	15'h4892: q<=8'hd8;
	15'h4893: q<=8'ha0;
	15'h4894: q<=8'hee;
	15'h4895: q<=8'ha2;
	15'h4896: q<=8'h1b;
	15'h4897: q<=8'h20;
	15'h4898: q<=8'ha9;
	15'h4899: q<=8'hd8;
	15'h489a: q<=8'ha5;
	15'h489b: q<=8'h09;
	15'h489c: q<=8'h4a;
	15'h489d: q<=8'h4a;
	15'h489e: q<=8'h4a;
	15'h489f: q<=8'h4a;
	15'h48a0: q<=8'h4a;
	15'h48a1: q<=8'haa;
	15'h48a2: q<=8'hbd;
	15'h48a3: q<=8'hc2;
	15'h48a4: q<=8'hd8;
	15'h48a5: q<=8'ha0;
	15'h48a6: q<=8'h32;
	15'h48a7: q<=8'ha2;
	15'h48a8: q<=8'hf8;
	15'h48a9: q<=8'h85;
	15'h48aa: q<=8'h29;
	15'h48ab: q<=8'h98;
	15'h48ac: q<=8'h20;
	15'h48ad: q<=8'h75;
	15'h48ae: q<=8'hdf;
	15'h48af: q<=8'ha9;
	15'h48b0: q<=8'h29;
	15'h48b1: q<=8'ha0;
	15'h48b2: q<=8'h01;
	15'h48b3: q<=8'h4c;
	15'h48b4: q<=8'hb1;
	15'h48b5: q<=8'hdf;
	15'h48b6: q<=8'h18;
	15'h48b7: q<=8'h18;
	15'h48b8: q<=8'h30;
	15'h48b9: q<=8'h50;
	15'h48ba: q<=8'h11;
	15'h48bb: q<=8'h14;
	15'h48bc: q<=8'h15;
	15'h48bd: q<=8'h16;
	15'h48be: q<=8'h21;
	15'h48bf: q<=8'h24;
	15'h48c0: q<=8'h25;
	15'h48c1: q<=8'h26;
	15'h48c2: q<=8'h00;
	15'h48c3: q<=8'h12;
	15'h48c4: q<=8'h14;
	15'h48c5: q<=8'h24;
	15'h48c6: q<=8'h15;
	15'h48c7: q<=8'h13;
	15'h48c8: q<=8'h00;
	15'h48c9: q<=8'h00;
	15'h48ca: q<=8'ha8;
	15'h48cb: q<=8'ha9;
	15'h48cc: q<=8'h00;
	15'h48cd: q<=8'h84;
	15'h48ce: q<=8'h79;
	15'h48cf: q<=8'h4a;
	15'h48d0: q<=8'h4a;
	15'h48d1: q<=8'h0a;
	15'h48d2: q<=8'haa;
	15'h48d3: q<=8'h98;
	15'h48d4: q<=8'h29;
	15'h48d5: q<=8'h0f;
	15'h48d6: q<=8'hd0;
	15'h48d7: q<=8'h01;
	15'h48d8: q<=8'he8;
	15'h48d9: q<=8'h9a;
	15'h48da: q<=8'ha9;
	15'h48db: q<=8'ha2;
	15'h48dc: q<=8'h8d;
	15'h48dd: q<=8'hc1;
	15'h48de: q<=8'h60;
	15'h48df: q<=8'hba;
	15'h48e0: q<=8'hd0;
	15'h48e1: q<=8'h07;
	15'h48e2: q<=8'ha9;
	15'h48e3: q<=8'h60;
	15'h48e4: q<=8'ha0;
	15'h48e5: q<=8'h09;
	15'h48e6: q<=8'hb8;
	15'h48e7: q<=8'h50;
	15'h48e8: q<=8'h04;
	15'h48e9: q<=8'ha9;
	15'h48ea: q<=8'hc0;
	15'h48eb: q<=8'ha0;
	15'h48ec: q<=8'h01;
	15'h48ed: q<=8'h8d;
	15'h48ee: q<=8'hc0;
	15'h48ef: q<=8'h60;
	15'h48f0: q<=8'ha9;
	15'h48f1: q<=8'h03;
	15'h48f2: q<=8'h8d;
	15'h48f3: q<=8'he0;
	15'h48f4: q<=8'h60;
	15'h48f5: q<=8'ha2;
	15'h48f6: q<=8'h00;
	15'h48f7: q<=8'h2c;
	15'h48f8: q<=8'h00;
	15'h48f9: q<=8'h0c;
	15'h48fa: q<=8'h30;
	15'h48fb: q<=8'hfb;
	15'h48fc: q<=8'h2c;
	15'h48fd: q<=8'h00;
	15'h48fe: q<=8'h0c;
	15'h48ff: q<=8'h10;
	15'h4900: q<=8'hfb;
	15'h4901: q<=8'h8d;
	15'h4902: q<=8'h00;
	15'h4903: q<=8'h50;
	15'h4904: q<=8'hca;
	15'h4905: q<=8'hd0;
	15'h4906: q<=8'hf0;
	15'h4907: q<=8'h88;
	15'h4908: q<=8'hd0;
	15'h4909: q<=8'hed;
	15'h490a: q<=8'h8e;
	15'h490b: q<=8'hc1;
	15'h490c: q<=8'h60;
	15'h490d: q<=8'ha9;
	15'h490e: q<=8'h00;
	15'h490f: q<=8'h8d;
	15'h4910: q<=8'he0;
	15'h4911: q<=8'h60;
	15'h4912: q<=8'ha0;
	15'h4913: q<=8'h09;
	15'h4914: q<=8'h2c;
	15'h4915: q<=8'h00;
	15'h4916: q<=8'h0c;
	15'h4917: q<=8'h30;
	15'h4918: q<=8'hfb;
	15'h4919: q<=8'h2c;
	15'h491a: q<=8'h00;
	15'h491b: q<=8'h0c;
	15'h491c: q<=8'h10;
	15'h491d: q<=8'hfb;
	15'h491e: q<=8'h8d;
	15'h491f: q<=8'h00;
	15'h4920: q<=8'h50;
	15'h4921: q<=8'hca;
	15'h4922: q<=8'hd0;
	15'h4923: q<=8'hf0;
	15'h4924: q<=8'h88;
	15'h4925: q<=8'hd0;
	15'h4926: q<=8'hed;
	15'h4927: q<=8'hba;
	15'h4928: q<=8'hca;
	15'h4929: q<=8'h9a;
	15'h492a: q<=8'h10;
	15'h492b: q<=8'hae;
	15'h492c: q<=8'h4c;
	15'h492d: q<=8'h0a;
	15'h492e: q<=8'hda;
	15'h492f: q<=8'h51;
	15'h4930: q<=8'h00;
	15'h4931: q<=8'ha8;
	15'h4932: q<=8'ha5;
	15'h4933: q<=8'h01;
	15'h4934: q<=8'hc9;
	15'h4935: q<=8'h20;
	15'h4936: q<=8'h90;
	15'h4937: q<=8'h02;
	15'h4938: q<=8'he9;
	15'h4939: q<=8'h18;
	15'h493a: q<=8'h29;
	15'h493b: q<=8'h1f;
	15'h493c: q<=8'h4c;
	15'h493d: q<=8'hcd;
	15'h493e: q<=8'hd8;
	15'h493f: q<=8'h78;
	15'h4940: q<=8'h8d;
	15'h4941: q<=8'h00;
	15'h4942: q<=8'h50;
	15'h4943: q<=8'h8d;
	15'h4944: q<=8'h00;
	15'h4945: q<=8'h58;
	15'h4946: q<=8'ha2;
	15'h4947: q<=8'hff;
	15'h4948: q<=8'h9a;
	15'h4949: q<=8'hd8;
	15'h494a: q<=8'he8;
	15'h494b: q<=8'h8a;
	15'h494c: q<=8'ha8;
	15'h494d: q<=8'h84;
	15'h494e: q<=8'h00;
	15'h494f: q<=8'h86;
	15'h4950: q<=8'h01;
	15'h4951: q<=8'ha0;
	15'h4952: q<=8'h00;
	15'h4953: q<=8'h91;
	15'h4954: q<=8'h00;
	15'h4955: q<=8'hc8;
	15'h4956: q<=8'hd0;
	15'h4957: q<=8'hfb;
	15'h4958: q<=8'he8;
	15'h4959: q<=8'he0;
	15'h495a: q<=8'h08;
	15'h495b: q<=8'hd0;
	15'h495c: q<=8'h02;
	15'h495d: q<=8'ha2;
	15'h495e: q<=8'h20;
	15'h495f: q<=8'he0;
	15'h4960: q<=8'h30;
	15'h4961: q<=8'h8d;
	15'h4962: q<=8'h00;
	15'h4963: q<=8'h50;
	15'h4964: q<=8'h90;
	15'h4965: q<=8'he7;
	15'h4966: q<=8'h85;
	15'h4967: q<=8'h01;
	15'h4968: q<=8'h8d;
	15'h4969: q<=8'he0;
	15'h496a: q<=8'h60;
	15'h496b: q<=8'h8d;
	15'h496c: q<=8'hcf;
	15'h496d: q<=8'h60;
	15'h496e: q<=8'h8d;
	15'h496f: q<=8'hdf;
	15'h4970: q<=8'h60;
	15'h4971: q<=8'ha2;
	15'h4972: q<=8'h07;
	15'h4973: q<=8'h8e;
	15'h4974: q<=8'hcf;
	15'h4975: q<=8'h60;
	15'h4976: q<=8'h8e;
	15'h4977: q<=8'hdf;
	15'h4978: q<=8'h60;
	15'h4979: q<=8'he8;
	15'h497a: q<=8'h9d;
	15'h497b: q<=8'hc0;
	15'h497c: q<=8'h60;
	15'h497d: q<=8'h9d;
	15'h497e: q<=8'hd0;
	15'h497f: q<=8'h60;
	15'h4980: q<=8'hca;
	15'h4981: q<=8'h10;
	15'h4982: q<=8'hf7;
	15'h4983: q<=8'had;
	15'h4984: q<=8'h00;
	15'h4985: q<=8'h0c;
	15'h4986: q<=8'h29;
	15'h4987: q<=8'h10;
	15'h4988: q<=8'hf0;
	15'h4989: q<=8'h1f;
	15'h498a: q<=8'h8d;
	15'h498b: q<=8'h00;
	15'h498c: q<=8'h50;
	15'h498d: q<=8'hce;
	15'h498e: q<=8'h00;
	15'h498f: q<=8'h01;
	15'h4990: q<=8'hd0;
	15'h4991: q<=8'hf8;
	15'h4992: q<=8'hce;
	15'h4993: q<=8'h01;
	15'h4994: q<=8'h01;
	15'h4995: q<=8'hd0;
	15'h4996: q<=8'hf3;
	15'h4997: q<=8'ha9;
	15'h4998: q<=8'h10;
	15'h4999: q<=8'h85;
	15'h499a: q<=8'hb4;
	15'h499b: q<=8'h20;
	15'h499c: q<=8'h11;
	15'h499d: q<=8'hde;
	15'h499e: q<=8'h20;
	15'h499f: q<=8'hac;
	15'h49a0: q<=8'hab;
	15'h49a1: q<=8'h20;
	15'h49a2: q<=8'h6e;
	15'h49a3: q<=8'hc1;
	15'h49a4: q<=8'h58;
	15'h49a5: q<=8'h4c;
	15'h49a6: q<=8'ha0;
	15'h49a7: q<=8'hc7;
	15'h49a8: q<=8'ha0;
	15'h49a9: q<=8'ha2;
	15'h49aa: q<=8'h11;
	15'h49ab: q<=8'h9a;
	15'h49ac: q<=8'ha0;
	15'h49ad: q<=8'h00;
	15'h49ae: q<=8'hba;
	15'h49af: q<=8'h96;
	15'h49b0: q<=8'h00;
	15'h49b1: q<=8'ha2;
	15'h49b2: q<=8'h01;
	15'h49b3: q<=8'hc8;
	15'h49b4: q<=8'hb9;
	15'h49b5: q<=8'h00;
	15'h49b6: q<=8'h00;
	15'h49b7: q<=8'hf0;
	15'h49b8: q<=8'h03;
	15'h49b9: q<=8'h4c;
	15'h49ba: q<=8'hca;
	15'h49bb: q<=8'hd8;
	15'h49bc: q<=8'he8;
	15'h49bd: q<=8'hd0;
	15'h49be: q<=8'hf4;
	15'h49bf: q<=8'hba;
	15'h49c0: q<=8'h8a;
	15'h49c1: q<=8'h8d;
	15'h49c2: q<=8'h00;
	15'h49c3: q<=8'h50;
	15'h49c4: q<=8'hc8;
	15'h49c5: q<=8'h59;
	15'h49c6: q<=8'h00;
	15'h49c7: q<=8'h00;
	15'h49c8: q<=8'hd0;
	15'h49c9: q<=8'hef;
	15'h49ca: q<=8'h99;
	15'h49cb: q<=8'h00;
	15'h49cc: q<=8'h00;
	15'h49cd: q<=8'hc8;
	15'h49ce: q<=8'hd0;
	15'h49cf: q<=8'hde;
	15'h49d0: q<=8'hba;
	15'h49d1: q<=8'h8a;
	15'h49d2: q<=8'h0a;
	15'h49d3: q<=8'haa;
	15'h49d4: q<=8'h90;
	15'h49d5: q<=8'hd5;
	15'h49d6: q<=8'ha0;
	15'h49d7: q<=8'h00;
	15'h49d8: q<=8'ha2;
	15'h49d9: q<=8'h01;
	15'h49da: q<=8'h84;
	15'h49db: q<=8'h00;
	15'h49dc: q<=8'h86;
	15'h49dd: q<=8'h01;
	15'h49de: q<=8'ha0;
	15'h49df: q<=8'h00;
	15'h49e0: q<=8'hb1;
	15'h49e1: q<=8'h00;
	15'h49e2: q<=8'hf0;
	15'h49e3: q<=8'h03;
	15'h49e4: q<=8'h4c;
	15'h49e5: q<=8'h31;
	15'h49e6: q<=8'hd9;
	15'h49e7: q<=8'ha9;
	15'h49e8: q<=8'h11;
	15'h49e9: q<=8'h91;
	15'h49ea: q<=8'h00;
	15'h49eb: q<=8'hd1;
	15'h49ec: q<=8'h00;
	15'h49ed: q<=8'hf0;
	15'h49ee: q<=8'h03;
	15'h49ef: q<=8'h4c;
	15'h49f0: q<=8'h2f;
	15'h49f1: q<=8'hd9;
	15'h49f2: q<=8'h0a;
	15'h49f3: q<=8'h90;
	15'h49f4: q<=8'hf4;
	15'h49f5: q<=8'ha9;
	15'h49f6: q<=8'h00;
	15'h49f7: q<=8'h91;
	15'h49f8: q<=8'h00;
	15'h49f9: q<=8'hc8;
	15'h49fa: q<=8'hd0;
	15'h49fb: q<=8'he4;
	15'h49fc: q<=8'h8d;
	15'h49fd: q<=8'h00;
	15'h49fe: q<=8'h50;
	15'h49ff: q<=8'he8;
	15'h4a00: q<=8'he0;
	15'h4a01: q<=8'h08;
	15'h4a02: q<=8'hd0;
	15'h4a03: q<=8'h02;
	15'h4a04: q<=8'ha2;
	15'h4a05: q<=8'h20;
	15'h4a06: q<=8'he0;
	15'h4a07: q<=8'h30;
	15'h4a08: q<=8'h90;
	15'h4a09: q<=8'hd0;
	15'h4a0a: q<=8'ha9;
	15'h4a0b: q<=8'h00;
	15'h4a0c: q<=8'ha8;
	15'h4a0d: q<=8'haa;
	15'h4a0e: q<=8'h85;
	15'h4a0f: q<=8'h3b;
	15'h4a10: q<=8'ha9;
	15'h4a11: q<=8'h30;
	15'h4a12: q<=8'h85;
	15'h4a13: q<=8'h3c;
	15'h4a14: q<=8'ha9;
	15'h4a15: q<=8'h08;
	15'h4a16: q<=8'h85;
	15'h4a17: q<=8'h38;
	15'h4a18: q<=8'h8a;
	15'h4a19: q<=8'h51;
	15'h4a1a: q<=8'h3b;
	15'h4a1b: q<=8'hc8;
	15'h4a1c: q<=8'hd0;
	15'h4a1d: q<=8'hfb;
	15'h4a1e: q<=8'he6;
	15'h4a1f: q<=8'h3c;
	15'h4a20: q<=8'h8d;
	15'h4a21: q<=8'h00;
	15'h4a22: q<=8'h50;
	15'h4a23: q<=8'hc6;
	15'h4a24: q<=8'h38;
	15'h4a25: q<=8'hd0;
	15'h4a26: q<=8'hf2;
	15'h4a27: q<=8'h95;
	15'h4a28: q<=8'h7d;
	15'h4a29: q<=8'he8;
	15'h4a2a: q<=8'he0;
	15'h4a2b: q<=8'h02;
	15'h4a2c: q<=8'hd0;
	15'h4a2d: q<=8'h04;
	15'h4a2e: q<=8'ha9;
	15'h4a2f: q<=8'h90;
	15'h4a30: q<=8'h85;
	15'h4a31: q<=8'h3c;
	15'h4a32: q<=8'he0;
	15'h4a33: q<=8'h0c;
	15'h4a34: q<=8'h90;
	15'h4a35: q<=8'hde;
	15'h4a36: q<=8'ha5;
	15'h4a37: q<=8'h7d;
	15'h4a38: q<=8'hf0;
	15'h4a39: q<=8'h0a;
	15'h4a3a: q<=8'ha9;
	15'h4a3b: q<=8'h40;
	15'h4a3c: q<=8'ha2;
	15'h4a3d: q<=8'ha4;
	15'h4a3e: q<=8'h8d;
	15'h4a3f: q<=8'hc4;
	15'h4a40: q<=8'h60;
	15'h4a41: q<=8'h8e;
	15'h4a42: q<=8'hc5;
	15'h4a43: q<=8'h60;
	15'h4a44: q<=8'ha2;
	15'h4a45: q<=8'h05;
	15'h4a46: q<=8'had;
	15'h4a47: q<=8'hca;
	15'h4a48: q<=8'h60;
	15'h4a49: q<=8'hcd;
	15'h4a4a: q<=8'hca;
	15'h4a4b: q<=8'h60;
	15'h4a4c: q<=8'hd0;
	15'h4a4d: q<=8'h05;
	15'h4a4e: q<=8'hca;
	15'h4a4f: q<=8'h10;
	15'h4a50: q<=8'hf8;
	15'h4a51: q<=8'h85;
	15'h4a52: q<=8'h7a;
	15'h4a53: q<=8'ha2;
	15'h4a54: q<=8'h05;
	15'h4a55: q<=8'had;
	15'h4a56: q<=8'hda;
	15'h4a57: q<=8'h60;
	15'h4a58: q<=8'hcd;
	15'h4a59: q<=8'hda;
	15'h4a5a: q<=8'h60;
	15'h4a5b: q<=8'hd0;
	15'h4a5c: q<=8'h05;
	15'h4a5d: q<=8'hca;
	15'h4a5e: q<=8'h10;
	15'h4a5f: q<=8'hf8;
	15'h4a60: q<=8'h85;
	15'h4a61: q<=8'h7b;
	15'h4a62: q<=8'h20;
	15'h4a63: q<=8'h11;
	15'h4a64: q<=8'hde;
	15'h4a65: q<=8'ha0;
	15'h4a66: q<=8'h02;
	15'h4a67: q<=8'had;
	15'h4a68: q<=8'hc9;
	15'h4a69: q<=8'h01;
	15'h4a6a: q<=8'hf0;
	15'h4a6b: q<=8'h0a;
	15'h4a6c: q<=8'h85;
	15'h4a6d: q<=8'h7c;
	15'h4a6e: q<=8'h20;
	15'h4a6f: q<=8'hf1;
	15'h4a70: q<=8'hdd;
	15'h4a71: q<=8'ha0;
	15'h4a72: q<=8'h00;
	15'h4a73: q<=8'h8c;
	15'h4a74: q<=8'hc9;
	15'h4a75: q<=8'h01;
	15'h4a76: q<=8'h84;
	15'h4a77: q<=8'h00;
	15'h4a78: q<=8'ha2;
	15'h4a79: q<=8'h07;
	15'h4a7a: q<=8'hbd;
	15'h4a7b: q<=8'hf9;
	15'h4a7c: q<=8'hda;
	15'h4a7d: q<=8'h9d;
	15'h4a7e: q<=8'h00;
	15'h4a7f: q<=8'h08;
	15'h4a80: q<=8'hca;
	15'h4a81: q<=8'h10;
	15'h4a82: q<=8'hf7;
	15'h4a83: q<=8'ha9;
	15'h4a84: q<=8'h00;
	15'h4a85: q<=8'h8d;
	15'h4a86: q<=8'he0;
	15'h4a87: q<=8'h60;
	15'h4a88: q<=8'ha9;
	15'h4a89: q<=8'h10;
	15'h4a8a: q<=8'h8d;
	15'h4a8b: q<=8'h00;
	15'h4a8c: q<=8'h40;
	15'h4a8d: q<=8'ha0;
	15'h4a8e: q<=8'h04;
	15'h4a8f: q<=8'ha2;
	15'h4a90: q<=8'h14;
	15'h4a91: q<=8'h2c;
	15'h4a92: q<=8'h00;
	15'h4a93: q<=8'h0c;
	15'h4a94: q<=8'h10;
	15'h4a95: q<=8'hfb;
	15'h4a96: q<=8'h2c;
	15'h4a97: q<=8'h00;
	15'h4a98: q<=8'h0c;
	15'h4a99: q<=8'h30;
	15'h4a9a: q<=8'hfb;
	15'h4a9b: q<=8'hca;
	15'h4a9c: q<=8'h10;
	15'h4a9d: q<=8'hf3;
	15'h4a9e: q<=8'h88;
	15'h4a9f: q<=8'h30;
	15'h4aa0: q<=8'h08;
	15'h4aa1: q<=8'h8d;
	15'h4aa2: q<=8'h00;
	15'h4aa3: q<=8'h50;
	15'h4aa4: q<=8'h2c;
	15'h4aa5: q<=8'h00;
	15'h4aa6: q<=8'h0c;
	15'h4aa7: q<=8'h50;
	15'h4aa8: q<=8'he6;
	15'h4aa9: q<=8'h8d;
	15'h4aaa: q<=8'h00;
	15'h4aab: q<=8'h58;
	15'h4aac: q<=8'ha9;
	15'h4aad: q<=8'h00;
	15'h4aae: q<=8'h85;
	15'h4aaf: q<=8'h74;
	15'h4ab0: q<=8'ha9;
	15'h4ab1: q<=8'h20;
	15'h4ab2: q<=8'h85;
	15'h4ab3: q<=8'h75;
	15'h4ab4: q<=8'h8d;
	15'h4ab5: q<=8'hcb;
	15'h4ab6: q<=8'h60;
	15'h4ab7: q<=8'had;
	15'h4ab8: q<=8'hc8;
	15'h4ab9: q<=8'h60;
	15'h4aba: q<=8'h85;
	15'h4abb: q<=8'h52;
	15'h4abc: q<=8'h29;
	15'h4abd: q<=8'h0f;
	15'h4abe: q<=8'h85;
	15'h4abf: q<=8'h50;
	15'h4ac0: q<=8'had;
	15'h4ac1: q<=8'h00;
	15'h4ac2: q<=8'h0c;
	15'h4ac3: q<=8'h49;
	15'h4ac4: q<=8'hff;
	15'h4ac5: q<=8'h29;
	15'h4ac6: q<=8'h2f;
	15'h4ac7: q<=8'h85;
	15'h4ac8: q<=8'h4e;
	15'h4ac9: q<=8'h29;
	15'h4aca: q<=8'h28;
	15'h4acb: q<=8'hf0;
	15'h4acc: q<=8'h0b;
	15'h4acd: q<=8'h06;
	15'h4ace: q<=8'h4c;
	15'h4acf: q<=8'h90;
	15'h4ad0: q<=8'h04;
	15'h4ad1: q<=8'he6;
	15'h4ad2: q<=8'h00;
	15'h4ad3: q<=8'he6;
	15'h4ad4: q<=8'h00;
	15'h4ad5: q<=8'hb8;
	15'h4ad6: q<=8'h50;
	15'h4ad7: q<=8'h04;
	15'h4ad8: q<=8'ha9;
	15'h4ad9: q<=8'h20;
	15'h4ada: q<=8'h85;
	15'h4adb: q<=8'h4c;
	15'h4adc: q<=8'h20;
	15'h4add: q<=8'h0f;
	15'h4ade: q<=8'hdb;
	15'h4adf: q<=8'h20;
	15'h4ae0: q<=8'h0d;
	15'h4ae1: q<=8'hdf;
	15'h4ae2: q<=8'h8d;
	15'h4ae3: q<=8'h00;
	15'h4ae4: q<=8'h48;
	15'h4ae5: q<=8'he6;
	15'h4ae6: q<=8'h03;
	15'h4ae7: q<=8'ha5;
	15'h4ae8: q<=8'h03;
	15'h4ae9: q<=8'h29;
	15'h4aea: q<=8'h03;
	15'h4aeb: q<=8'hd0;
	15'h4aec: q<=8'h03;
	15'h4aed: q<=8'h20;
	15'h4aee: q<=8'h1b;
	15'h4aef: q<=8'hde;
	15'h4af0: q<=8'had;
	15'h4af1: q<=8'h00;
	15'h4af2: q<=8'h0c;
	15'h4af3: q<=8'h29;
	15'h4af4: q<=8'h10;
	15'h4af5: q<=8'hf0;
	15'h4af6: q<=8'h96;
	15'h4af7: q<=8'hd0;
	15'h4af8: q<=8'hfe;
	15'h4af9: q<=8'h00;
	15'h4afa: q<=8'h04;
	15'h4afb: q<=8'h08;
	15'h4afc: q<=8'h0c;
	15'h4afd: q<=8'h03;
	15'h4afe: q<=8'h07;
	15'h4aff: q<=8'h0b;
	15'h4b00: q<=8'h0b;
	15'h4b01: q<=8'h59;
	15'h4b02: q<=8'hdb;
	15'h4b03: q<=8'hf6;
	15'h4b04: q<=8'hdb;
	15'h4b05: q<=8'h83;
	15'h4b06: q<=8'hdb;
	15'h4b07: q<=8'h99;
	15'h4b08: q<=8'hdb;
	15'h4b09: q<=8'h7d;
	15'h4b0a: q<=8'hdb;
	15'h4b0b: q<=8'h6e;
	15'h4b0c: q<=8'hdb;
	15'h4b0d: q<=8'h21;
	15'h4b0e: q<=8'hdb;
	15'h4b0f: q<=8'ha6;
	15'h4b10: q<=8'h00;
	15'h4b11: q<=8'he0;
	15'h4b12: q<=8'h0e;
	15'h4b13: q<=8'h90;
	15'h4b14: q<=8'h04;
	15'h4b15: q<=8'ha2;
	15'h4b16: q<=8'h02;
	15'h4b17: q<=8'h86;
	15'h4b18: q<=8'h00;
	15'h4b19: q<=8'hbd;
	15'h4b1a: q<=8'h02;
	15'h4b1b: q<=8'hdb;
	15'h4b1c: q<=8'h48;
	15'h4b1d: q<=8'hbd;
	15'h4b1e: q<=8'h01;
	15'h4b1f: q<=8'hdb;
	15'h4b20: q<=8'h48;
	15'h4b21: q<=8'h60;
	15'h4b22: q<=8'ha9;
	15'h4b23: q<=8'h00;
	15'h4b24: q<=8'h8d;
	15'h4b25: q<=8'he0;
	15'h4b26: q<=8'h60;
	15'h4b27: q<=8'h8d;
	15'h4b28: q<=8'h80;
	15'h4b29: q<=8'h60;
	15'h4b2a: q<=8'h8d;
	15'h4b2b: q<=8'hc0;
	15'h4b2c: q<=8'h60;
	15'h4b2d: q<=8'h8d;
	15'h4b2e: q<=8'hd0;
	15'h4b2f: q<=8'h60;
	15'h4b30: q<=8'h8d;
	15'h4b31: q<=8'h00;
	15'h4b32: q<=8'h60;
	15'h4b33: q<=8'h8d;
	15'h4b34: q<=8'h40;
	15'h4b35: q<=8'h60;
	15'h4b36: q<=8'had;
	15'h4b37: q<=8'h40;
	15'h4b38: q<=8'h60;
	15'h4b39: q<=8'had;
	15'h4b3a: q<=8'h60;
	15'h4b3b: q<=8'h60;
	15'h4b3c: q<=8'had;
	15'h4b3d: q<=8'h70;
	15'h4b3e: q<=8'h60;
	15'h4b3f: q<=8'had;
	15'h4b40: q<=8'h50;
	15'h4b41: q<=8'h60;
	15'h4b42: q<=8'ha9;
	15'h4b43: q<=8'h08;
	15'h4b44: q<=8'h8d;
	15'h4b45: q<=8'he0;
	15'h4b46: q<=8'h60;
	15'h4b47: q<=8'ha9;
	15'h4b48: q<=8'h01;
	15'h4b49: q<=8'ha2;
	15'h4b4a: q<=8'h1f;
	15'h4b4b: q<=8'h18;
	15'h4b4c: q<=8'h9d;
	15'h4b4d: q<=8'h80;
	15'h4b4e: q<=8'h60;
	15'h4b4f: q<=8'h2a;
	15'h4b50: q<=8'hca;
	15'h4b51: q<=8'h10;
	15'h4b52: q<=8'hf9;
	15'h4b53: q<=8'ha9;
	15'h4b54: q<=8'h34;
	15'h4b55: q<=8'ha2;
	15'h4b56: q<=8'ha6;
	15'h4b57: q<=8'h4c;
	15'h4b58: q<=8'h39;
	15'h4b59: q<=8'hdf;
	15'h4b5a: q<=8'had;
	15'h4b5b: q<=8'hca;
	15'h4b5c: q<=8'h01;
	15'h4b5d: q<=8'h0d;
	15'h4b5e: q<=8'hc7;
	15'h4b5f: q<=8'h01;
	15'h4b60: q<=8'hd0;
	15'h4b61: q<=8'h0c;
	15'h4b62: q<=8'h20;
	15'h4b63: q<=8'h11;
	15'h4b64: q<=8'hde;
	15'h4b65: q<=8'had;
	15'h4b66: q<=8'hc9;
	15'h4b67: q<=8'h01;
	15'h4b68: q<=8'h85;
	15'h4b69: q<=8'h7c;
	15'h4b6a: q<=8'ha9;
	15'h4b6b: q<=8'h02;
	15'h4b6c: q<=8'h85;
	15'h4b6d: q<=8'h00;
	15'h4b6e: q<=8'h60;
	15'h4b6f: q<=8'ha5;
	15'h4b70: q<=8'h50;
	15'h4b71: q<=8'h4a;
	15'h4b72: q<=8'ha8;
	15'h4b73: q<=8'ha9;
	15'h4b74: q<=8'h68;
	15'h4b75: q<=8'h20;
	15'h4b76: q<=8'h4c;
	15'h4b77: q<=8'hdf;
	15'h4b78: q<=8'ha2;
	15'h4b79: q<=8'h4e;
	15'h4b7a: q<=8'ha9;
	15'h4b7b: q<=8'h33;
	15'h4b7c: q<=8'hd0;
	15'h4b7d: q<=8'h0a;
	15'h4b7e: q<=8'ha2;
	15'h4b7f: q<=8'hb6;
	15'h4b80: q<=8'ha9;
	15'h4b81: q<=8'h32;
	15'h4b82: q<=8'hd0;
	15'h4b83: q<=8'h04;
	15'h4b84: q<=8'ha9;
	15'h4b85: q<=8'h33;
	15'h4b86: q<=8'ha2;
	15'h4b87: q<=8'h0a;
	15'h4b88: q<=8'h20;
	15'h4b89: q<=8'h39;
	15'h4b8a: q<=8'hdf;
	15'h4b8b: q<=8'ha2;
	15'h4b8c: q<=8'h06;
	15'h4b8d: q<=8'ha9;
	15'h4b8e: q<=8'h00;
	15'h4b8f: q<=8'h9d;
	15'h4b90: q<=8'hc1;
	15'h4b91: q<=8'h60;
	15'h4b92: q<=8'h9d;
	15'h4b93: q<=8'hd1;
	15'h4b94: q<=8'h60;
	15'h4b95: q<=8'hca;
	15'h4b96: q<=8'hca;
	15'h4b97: q<=8'h10;
	15'h4b98: q<=8'hf6;
	15'h4b99: q<=8'h60;
	15'h4b9a: q<=8'ha5;
	15'h4b9b: q<=8'h03;
	15'h4b9c: q<=8'h29;
	15'h4b9d: q<=8'h3f;
	15'h4b9e: q<=8'hd0;
	15'h4b9f: q<=8'h02;
	15'h4ba0: q<=8'he6;
	15'h4ba1: q<=8'h39;
	15'h4ba2: q<=8'ha5;
	15'h4ba3: q<=8'h39;
	15'h4ba4: q<=8'h29;
	15'h4ba5: q<=8'h07;
	15'h4ba6: q<=8'haa;
	15'h4ba7: q<=8'hbc;
	15'h4ba8: q<=8'hd5;
	15'h4ba9: q<=8'hdb;
	15'h4baa: q<=8'ha9;
	15'h4bab: q<=8'h00;
	15'h4bac: q<=8'h99;
	15'h4bad: q<=8'hc1;
	15'h4bae: q<=8'h60;
	15'h4baf: q<=8'hbc;
	15'h4bb0: q<=8'hd6;
	15'h4bb1: q<=8'hdb;
	15'h4bb2: q<=8'hbd;
	15'h4bb3: q<=8'hdc;
	15'h4bb4: q<=8'hdf;
	15'h4bb5: q<=8'h99;
	15'h4bb6: q<=8'hc0;
	15'h4bb7: q<=8'h60;
	15'h4bb8: q<=8'ha9;
	15'h4bb9: q<=8'ha8;
	15'h4bba: q<=8'h99;
	15'h4bbb: q<=8'hc1;
	15'h4bbc: q<=8'h60;
	15'h4bbd: q<=8'ha9;
	15'h4bbe: q<=8'h34;
	15'h4bbf: q<=8'ha2;
	15'h4bc0: q<=8'h56;
	15'h4bc1: q<=8'h20;
	15'h4bc2: q<=8'h39;
	15'h4bc3: q<=8'hdf;
	15'h4bc4: q<=8'ha5;
	15'h4bc5: q<=8'h03;
	15'h4bc6: q<=8'h29;
	15'h4bc7: q<=8'h7f;
	15'h4bc8: q<=8'ha8;
	15'h4bc9: q<=8'ha9;
	15'h4bca: q<=8'h01;
	15'h4bcb: q<=8'h20;
	15'h4bcc: q<=8'h6c;
	15'h4bcd: q<=8'hdf;
	15'h4bce: q<=8'ha9;
	15'h4bcf: q<=8'h34;
	15'h4bd0: q<=8'ha2;
	15'h4bd1: q<=8'haa;
	15'h4bd2: q<=8'h4c;
	15'h4bd3: q<=8'h39;
	15'h4bd4: q<=8'hdf;
	15'h4bd5: q<=8'h16;
	15'h4bd6: q<=8'h00;
	15'h4bd7: q<=8'h10;
	15'h4bd8: q<=8'h02;
	15'h4bd9: q<=8'h12;
	15'h4bda: q<=8'h04;
	15'h4bdb: q<=8'h14;
	15'h4bdc: q<=8'h06;
	15'h4bdd: q<=8'h16;
	15'h4bde: q<=8'h00;
	15'h4bdf: q<=8'hea;
	15'h4be0: q<=8'h8d;
	15'h4be1: q<=8'hdb;
	15'h4be2: q<=8'h60;
	15'h4be3: q<=8'had;
	15'h4be4: q<=8'hd8;
	15'h4be5: q<=8'h60;
	15'h4be6: q<=8'h29;
	15'h4be7: q<=8'h07;
	15'h4be8: q<=8'h85;
	15'h4be9: q<=8'h37;
	15'h4bea: q<=8'h8d;
	15'h4beb: q<=8'hcb;
	15'h4bec: q<=8'h60;
	15'h4bed: q<=8'had;
	15'h4bee: q<=8'hc8;
	15'h4bef: q<=8'h60;
	15'h4bf0: q<=8'h29;
	15'h4bf1: q<=8'h20;
	15'h4bf2: q<=8'h4a;
	15'h4bf3: q<=8'h4a;
	15'h4bf4: q<=8'h05;
	15'h4bf5: q<=8'h37;
	15'h4bf6: q<=8'h60;
	15'h4bf7: q<=8'ha5;
	15'h4bf8: q<=8'h2e;
	15'h4bf9: q<=8'hf0;
	15'h4bfa: q<=8'h1e;
	15'h4bfb: q<=8'h8d;
	15'h4bfc: q<=8'h95;
	15'h4bfd: q<=8'h60;
	15'h4bfe: q<=8'h8d;
	15'h4bff: q<=8'h8d;
	15'h4c00: q<=8'h60;
	15'h4c01: q<=8'ha5;
	15'h4c02: q<=8'h2f;
	15'h4c03: q<=8'h8d;
	15'h4c04: q<=8'h96;
	15'h4c05: q<=8'h60;
	15'h4c06: q<=8'ha2;
	15'h4c07: q<=8'h00;
	15'h4c08: q<=8'h20;
	15'h4c09: q<=8'he6;
	15'h4c0a: q<=8'hdc;
	15'h4c0b: q<=8'hc9;
	15'h4c0c: q<=8'h01;
	15'h4c0d: q<=8'hd0;
	15'h4c0e: q<=8'h06;
	15'h4c0f: q<=8'h98;
	15'h4c10: q<=8'hd0;
	15'h4c11: q<=8'h03;
	15'h4c12: q<=8'h8a;
	15'h4c13: q<=8'h10;
	15'h4c14: q<=8'h04;
	15'h4c15: q<=8'ha9;
	15'h4c16: q<=8'hff;
	15'h4c17: q<=8'h85;
	15'h4c18: q<=8'h78;
	15'h4c19: q<=8'ha2;
	15'h4c1a: q<=8'h00;
	15'h4c1b: q<=8'h86;
	15'h4c1c: q<=8'h73;
	15'h4c1d: q<=8'he6;
	15'h4c1e: q<=8'h2e;
	15'h4c1f: q<=8'hd0;
	15'h4c20: q<=8'h06;
	15'h4c21: q<=8'he6;
	15'h4c22: q<=8'h2f;
	15'h4c23: q<=8'h10;
	15'h4c24: q<=8'h02;
	15'h4c25: q<=8'h86;
	15'h4c26: q<=8'h2f;
	15'h4c27: q<=8'h8d;
	15'h4c28: q<=8'hdb;
	15'h4c29: q<=8'h60;
	15'h4c2a: q<=8'had;
	15'h4c2b: q<=8'hd8;
	15'h4c2c: q<=8'h60;
	15'h4c2d: q<=8'h29;
	15'h4c2e: q<=8'h78;
	15'h4c2f: q<=8'h85;
	15'h4c30: q<=8'h4d;
	15'h4c31: q<=8'hf0;
	15'h4c32: q<=8'h05;
	15'h4c33: q<=8'h8d;
	15'h4c34: q<=8'hc0;
	15'h4c35: q<=8'h60;
	15'h4c36: q<=8'ha2;
	15'h4c37: q<=8'ha4;
	15'h4c38: q<=8'h8e;
	15'h4c39: q<=8'hc1;
	15'h4c3a: q<=8'h60;
	15'h4c3b: q<=8'ha2;
	15'h4c3c: q<=8'h00;
	15'h4c3d: q<=8'ha5;
	15'h4c3e: q<=8'h4e;
	15'h4c3f: q<=8'hf0;
	15'h4c40: q<=8'h06;
	15'h4c41: q<=8'h0a;
	15'h4c42: q<=8'h8d;
	15'h4c43: q<=8'hc2;
	15'h4c44: q<=8'h60;
	15'h4c45: q<=8'ha2;
	15'h4c46: q<=8'ha4;
	15'h4c47: q<=8'h8e;
	15'h4c48: q<=8'hc3;
	15'h4c49: q<=8'h60;
	15'h4c4a: q<=8'h20;
	15'h4c4b: q<=8'h0d;
	15'h4c4c: q<=8'hdd;
	15'h4c4d: q<=8'ha4;
	15'h4c4e: q<=8'h4d;
	15'h4c4f: q<=8'ha9;
	15'h4c50: q<=8'hd0;
	15'h4c51: q<=8'ha2;
	15'h4c52: q<=8'hf0;
	15'h4c53: q<=8'h20;
	15'h4c54: q<=8'h2b;
	15'h4c55: q<=8'hdd;
	15'h4c56: q<=8'ha4;
	15'h4c57: q<=8'h4e;
	15'h4c58: q<=8'h20;
	15'h4c59: q<=8'h27;
	15'h4c5a: q<=8'hdd;
	15'h4c5b: q<=8'ha5;
	15'h4c5c: q<=8'h52;
	15'h4c5d: q<=8'h29;
	15'h4c5e: q<=8'h10;
	15'h4c5f: q<=8'hf0;
	15'h4c60: q<=8'h1d;
	15'h4c61: q<=8'ha9;
	15'h4c62: q<=8'h34;
	15'h4c63: q<=8'ha2;
	15'h4c64: q<=8'h82;
	15'h4c65: q<=8'h20;
	15'h4c66: q<=8'h39;
	15'h4c67: q<=8'hdf;
	15'h4c68: q<=8'ha0;
	15'h4c69: q<=8'h10;
	15'h4c6a: q<=8'ha5;
	15'h4c6b: q<=8'h4d;
	15'h4c6c: q<=8'h29;
	15'h4c6d: q<=8'h60;
	15'h4c6e: q<=8'hf0;
	15'h4c6f: q<=8'h0e;
	15'h4c70: q<=8'h49;
	15'h4c71: q<=8'h20;
	15'h4c72: q<=8'hf0;
	15'h4c73: q<=8'h04;
	15'h4c74: q<=8'ha9;
	15'h4c75: q<=8'h04;
	15'h4c76: q<=8'ha0;
	15'h4c77: q<=8'h08;
	15'h4c78: q<=8'h8d;
	15'h4c79: q<=8'he0;
	15'h4c7a: q<=8'h60;
	15'h4c7b: q<=8'h8c;
	15'h4c7c: q<=8'h00;
	15'h4c7d: q<=8'h40;
	15'h4c7e: q<=8'ha9;
	15'h4c7f: q<=8'h34;
	15'h4c80: q<=8'ha2;
	15'h4c81: q<=8'h92;
	15'h4c82: q<=8'h20;
	15'h4c83: q<=8'h39;
	15'h4c84: q<=8'hdf;
	15'h4c85: q<=8'ha2;
	15'h4c86: q<=8'h0b;
	15'h4c87: q<=8'hb5;
	15'h4c88: q<=8'h7d;
	15'h4c89: q<=8'hf0;
	15'h4c8a: q<=8'h19;
	15'h4c8b: q<=8'h85;
	15'h4c8c: q<=8'h35;
	15'h4c8d: q<=8'h86;
	15'h4c8e: q<=8'h38;
	15'h4c8f: q<=8'h8a;
	15'h4c90: q<=8'h20;
	15'h4c91: q<=8'h1f;
	15'h4c92: q<=8'hdf;
	15'h4c93: q<=8'ha0;
	15'h4c94: q<=8'hf4;
	15'h4c95: q<=8'ha2;
	15'h4c96: q<=8'hf4;
	15'h4c97: q<=8'ha5;
	15'h4c98: q<=8'h35;
	15'h4c99: q<=8'h20;
	15'h4c9a: q<=8'ha9;
	15'h4c9b: q<=8'hd8;
	15'h4c9c: q<=8'ha9;
	15'h4c9d: q<=8'h0c;
	15'h4c9e: q<=8'haa;
	15'h4c9f: q<=8'h20;
	15'h4ca0: q<=8'h75;
	15'h4ca1: q<=8'hdf;
	15'h4ca2: q<=8'ha6;
	15'h4ca3: q<=8'h38;
	15'h4ca4: q<=8'hca;
	15'h4ca5: q<=8'h10;
	15'h4ca6: q<=8'he0;
	15'h4ca7: q<=8'h20;
	15'h4ca8: q<=8'h53;
	15'h4ca9: q<=8'hdf;
	15'h4caa: q<=8'ha9;
	15'h4cab: q<=8'h00;
	15'h4cac: q<=8'ha2;
	15'h4cad: q<=8'h16;
	15'h4cae: q<=8'h20;
	15'h4caf: q<=8'h75;
	15'h4cb0: q<=8'hdf;
	15'h4cb1: q<=8'ha2;
	15'h4cb2: q<=8'h04;
	15'h4cb3: q<=8'h86;
	15'h4cb4: q<=8'h37;
	15'h4cb5: q<=8'ha6;
	15'h4cb6: q<=8'h37;
	15'h4cb7: q<=8'ha0;
	15'h4cb8: q<=8'h00;
	15'h4cb9: q<=8'hb5;
	15'h4cba: q<=8'h78;
	15'h4cbb: q<=8'hf0;
	15'h4cbc: q<=8'h03;
	15'h4cbd: q<=8'hbc;
	15'h4cbe: q<=8'he1;
	15'h4cbf: q<=8'hdc;
	15'h4cc0: q<=8'hb9;
	15'h4cc1: q<=8'he4;
	15'h4cc2: q<=8'h31;
	15'h4cc3: q<=8'hbe;
	15'h4cc4: q<=8'he5;
	15'h4cc5: q<=8'h31;
	15'h4cc6: q<=8'h20;
	15'h4cc7: q<=8'h57;
	15'h4cc8: q<=8'hdf;
	15'h4cc9: q<=8'hc6;
	15'h4cca: q<=8'h37;
	15'h4ccb: q<=8'h10;
	15'h4ccc: q<=8'he8;
	15'h4ccd: q<=8'ha2;
	15'h4cce: q<=8'hac;
	15'h4ccf: q<=8'ha9;
	15'h4cd0: q<=8'h30;
	15'h4cd1: q<=8'h20;
	15'h4cd2: q<=8'h75;
	15'h4cd3: q<=8'hdf;
	15'h4cd4: q<=8'ha4;
	15'h4cd5: q<=8'h50;
	15'h4cd6: q<=8'hb9;
	15'h4cd7: q<=8'he8;
	15'h4cd8: q<=8'hdf;
	15'h4cd9: q<=8'hbe;
	15'h4cda: q<=8'he4;
	15'h4cdb: q<=8'hdf;
	15'h4cdc: q<=8'ha0;
	15'h4cdd: q<=8'hc0;
	15'h4cde: q<=8'h4c;
	15'h4cdf: q<=8'h73;
	15'h4ce0: q<=8'hdf;
	15'h4ce1: q<=8'h2e;
	15'h4ce2: q<=8'h38;
	15'h4ce3: q<=8'h34;
	15'h4ce4: q<=8'h36;
	15'h4ce5: q<=8'h1e;
	15'h4ce6: q<=8'ha0;
	15'h4ce7: q<=8'h00;
	15'h4ce8: q<=8'h84;
	15'h4ce9: q<=8'h73;
	15'h4cea: q<=8'h8c;
	15'h4ceb: q<=8'h14;
	15'h4cec: q<=8'h04;
	15'h4ced: q<=8'h8d;
	15'h4cee: q<=8'h8e;
	15'h4cef: q<=8'h60;
	15'h4cf0: q<=8'h8e;
	15'h4cf1: q<=8'h8f;
	15'h4cf2: q<=8'h60;
	15'h4cf3: q<=8'h8c;
	15'h4cf4: q<=8'h90;
	15'h4cf5: q<=8'h60;
	15'h4cf6: q<=8'ha2;
	15'h4cf7: q<=8'h10;
	15'h4cf8: q<=8'h8e;
	15'h4cf9: q<=8'h8c;
	15'h4cfa: q<=8'h60;
	15'h4cfb: q<=8'h8e;
	15'h4cfc: q<=8'h94;
	15'h4cfd: q<=8'h60;
	15'h4cfe: q<=8'hca;
	15'h4cff: q<=8'h30;
	15'h4d00: q<=8'h0b;
	15'h4d01: q<=8'had;
	15'h4d02: q<=8'h40;
	15'h4d03: q<=8'h60;
	15'h4d04: q<=8'h30;
	15'h4d05: q<=8'hf8;
	15'h4d06: q<=8'had;
	15'h4d07: q<=8'h60;
	15'h4d08: q<=8'h60;
	15'h4d09: q<=8'hac;
	15'h4d0a: q<=8'h70;
	15'h4d0b: q<=8'h60;
	15'h4d0c: q<=8'h60;
	15'h4d0d: q<=8'h20;
	15'h4d0e: q<=8'h53;
	15'h4d0f: q<=8'hdf;
	15'h4d10: q<=8'ha9;
	15'h4d11: q<=8'h00;
	15'h4d12: q<=8'h20;
	15'h4d13: q<=8'h6a;
	15'h4d14: q<=8'hdf;
	15'h4d15: q<=8'ha9;
	15'h4d16: q<=8'he8;
	15'h4d17: q<=8'hac;
	15'h4d18: q<=8'h00;
	15'h4d19: q<=8'h0d;
	15'h4d1a: q<=8'h20;
	15'h4d1b: q<=8'h29;
	15'h4d1c: q<=8'hdd;
	15'h4d1d: q<=8'hac;
	15'h4d1e: q<=8'h00;
	15'h4d1f: q<=8'h0e;
	15'h4d20: q<=8'h20;
	15'h4d21: q<=8'h27;
	15'h4d22: q<=8'hdd;
	15'h4d23: q<=8'h20;
	15'h4d24: q<=8'he0;
	15'h4d25: q<=8'hdb;
	15'h4d26: q<=8'ha8;
	15'h4d27: q<=8'ha9;
	15'h4d28: q<=8'hd0;
	15'h4d29: q<=8'ha2;
	15'h4d2a: q<=8'hf8;
	15'h4d2b: q<=8'h84;
	15'h4d2c: q<=8'h35;
	15'h4d2d: q<=8'h20;
	15'h4d2e: q<=8'h75;
	15'h4d2f: q<=8'hdf;
	15'h4d30: q<=8'ha2;
	15'h4d31: q<=8'h07;
	15'h4d32: q<=8'h86;
	15'h4d33: q<=8'h37;
	15'h4d34: q<=8'h06;
	15'h4d35: q<=8'h35;
	15'h4d36: q<=8'ha9;
	15'h4d37: q<=8'h00;
	15'h4d38: q<=8'h2a;
	15'h4d39: q<=8'h20;
	15'h4d3a: q<=8'h1f;
	15'h4d3b: q<=8'hdf;
	15'h4d3c: q<=8'hc6;
	15'h4d3d: q<=8'h37;
	15'h4d3e: q<=8'h10;
	15'h4d3f: q<=8'hf4;
	15'h4d40: q<=8'h60;
	15'h4d41: q<=8'had;
	15'h4d42: q<=8'h0f;
	15'h4d43: q<=8'h04;
	15'h4d44: q<=8'h0a;
	15'h4d45: q<=8'h85;
	15'h4d46: q<=8'h29;
	15'h4d47: q<=8'had;
	15'h4d48: q<=8'h10;
	15'h4d49: q<=8'h04;
	15'h4d4a: q<=8'h2a;
	15'h4d4b: q<=8'h85;
	15'h4d4c: q<=8'h2a;
	15'h4d4d: q<=8'had;
	15'h4d4e: q<=8'h0c;
	15'h4d4f: q<=8'h04;
	15'h4d50: q<=8'h18;
	15'h4d51: q<=8'h65;
	15'h4d52: q<=8'h29;
	15'h4d53: q<=8'h8d;
	15'h4d54: q<=8'h95;
	15'h4d55: q<=8'h60;
	15'h4d56: q<=8'h85;
	15'h4d57: q<=8'h29;
	15'h4d58: q<=8'had;
	15'h4d59: q<=8'h0d;
	15'h4d5a: q<=8'h04;
	15'h4d5b: q<=8'h65;
	15'h4d5c: q<=8'h2a;
	15'h4d5d: q<=8'h8d;
	15'h4d5e: q<=8'h96;
	15'h4d5f: q<=8'h60;
	15'h4d60: q<=8'h05;
	15'h4d61: q<=8'h29;
	15'h4d62: q<=8'hd0;
	15'h4d63: q<=8'h05;
	15'h4d64: q<=8'ha9;
	15'h4d65: q<=8'h01;
	15'h4d66: q<=8'h8d;
	15'h4d67: q<=8'h95;
	15'h4d68: q<=8'h60;
	15'h4d69: q<=8'had;
	15'h4d6a: q<=8'h09;
	15'h4d6b: q<=8'h04;
	15'h4d6c: q<=8'h8d;
	15'h4d6d: q<=8'h8d;
	15'h4d6e: q<=8'h60;
	15'h4d6f: q<=8'had;
	15'h4d70: q<=8'h0a;
	15'h4d71: q<=8'h04;
	15'h4d72: q<=8'hae;
	15'h4d73: q<=8'h0b;
	15'h4d74: q<=8'h04;
	15'h4d75: q<=8'h20;
	15'h4d76: q<=8'he6;
	15'h4d77: q<=8'hdc;
	15'h4d78: q<=8'h8d;
	15'h4d79: q<=8'h12;
	15'h4d7a: q<=8'h04;
	15'h4d7b: q<=8'h8c;
	15'h4d7c: q<=8'h13;
	15'h4d7d: q<=8'h04;
	15'h4d7e: q<=8'ha9;
	15'h4d7f: q<=8'h3d;
	15'h4d80: q<=8'ha2;
	15'h4d81: q<=8'hce;
	15'h4d82: q<=8'h20;
	15'h4d83: q<=8'h39;
	15'h4d84: q<=8'hdf;
	15'h4d85: q<=8'ha9;
	15'h4d86: q<=8'h06;
	15'h4d87: q<=8'h85;
	15'h4d88: q<=8'h3b;
	15'h4d89: q<=8'ha9;
	15'h4d8a: q<=8'h04;
	15'h4d8b: q<=8'h85;
	15'h4d8c: q<=8'h3c;
	15'h4d8d: q<=8'h85;
	15'h4d8e: q<=8'h37;
	15'h4d8f: q<=8'ha0;
	15'h4d90: q<=8'h00;
	15'h4d91: q<=8'h84;
	15'h4d92: q<=8'h31;
	15'h4d93: q<=8'h84;
	15'h4d94: q<=8'h32;
	15'h4d95: q<=8'h84;
	15'h4d96: q<=8'h33;
	15'h4d97: q<=8'h84;
	15'h4d98: q<=8'h34;
	15'h4d99: q<=8'hb1;
	15'h4d9a: q<=8'h3b;
	15'h4d9b: q<=8'h85;
	15'h4d9c: q<=8'h56;
	15'h4d9d: q<=8'he6;
	15'h4d9e: q<=8'h3b;
	15'h4d9f: q<=8'hb1;
	15'h4da0: q<=8'h3b;
	15'h4da1: q<=8'h85;
	15'h4da2: q<=8'h57;
	15'h4da3: q<=8'he6;
	15'h4da4: q<=8'h3b;
	15'h4da5: q<=8'hb1;
	15'h4da6: q<=8'h3b;
	15'h4da7: q<=8'h85;
	15'h4da8: q<=8'h58;
	15'h4da9: q<=8'he6;
	15'h4daa: q<=8'h3b;
	15'h4dab: q<=8'hf8;
	15'h4dac: q<=8'ha0;
	15'h4dad: q<=8'h17;
	15'h4dae: q<=8'h84;
	15'h4daf: q<=8'h38;
	15'h4db0: q<=8'h26;
	15'h4db1: q<=8'h56;
	15'h4db2: q<=8'h26;
	15'h4db3: q<=8'h57;
	15'h4db4: q<=8'h26;
	15'h4db5: q<=8'h58;
	15'h4db6: q<=8'ha0;
	15'h4db7: q<=8'h03;
	15'h4db8: q<=8'ha2;
	15'h4db9: q<=8'h00;
	15'h4dba: q<=8'hb5;
	15'h4dbb: q<=8'h31;
	15'h4dbc: q<=8'h75;
	15'h4dbd: q<=8'h31;
	15'h4dbe: q<=8'h95;
	15'h4dbf: q<=8'h31;
	15'h4dc0: q<=8'he8;
	15'h4dc1: q<=8'h88;
	15'h4dc2: q<=8'h10;
	15'h4dc3: q<=8'hf6;
	15'h4dc4: q<=8'hc6;
	15'h4dc5: q<=8'h38;
	15'h4dc6: q<=8'h10;
	15'h4dc7: q<=8'he8;
	15'h4dc8: q<=8'hd8;
	15'h4dc9: q<=8'ha9;
	15'h4dca: q<=8'h31;
	15'h4dcb: q<=8'ha0;
	15'h4dcc: q<=8'h04;
	15'h4dcd: q<=8'h20;
	15'h4dce: q<=8'hb1;
	15'h4dcf: q<=8'hdf;
	15'h4dd0: q<=8'ha9;
	15'h4dd1: q<=8'hd0;
	15'h4dd2: q<=8'ha2;
	15'h4dd3: q<=8'hf8;
	15'h4dd4: q<=8'h20;
	15'h4dd5: q<=8'h75;
	15'h4dd6: q<=8'hdf;
	15'h4dd7: q<=8'hc6;
	15'h4dd8: q<=8'h37;
	15'h4dd9: q<=8'h10;
	15'h4dda: q<=8'hb4;
	15'h4ddb: q<=8'h60;
	15'h4ddc: q<=8'h73;
	15'h4ddd: q<=8'h00;
	15'h4dde: q<=8'h09;
	15'h4ddf: q<=8'h0a;
	15'h4de0: q<=8'h15;
	15'h4de1: q<=8'h16;
	15'h4de2: q<=8'h22;
	15'h4de3: q<=8'h15;
	15'h4de4: q<=8'h06;
	15'h4de5: q<=8'h15;
	15'h4de6: q<=8'h07;
	15'h4de7: q<=8'h06;
	15'h4de8: q<=8'h04;
	15'h4de9: q<=8'ha9;
	15'h4dea: q<=8'h04;
	15'h4deb: q<=8'hd0;
	15'h4dec: q<=8'h06;
	15'h4ded: q<=8'ha9;
	15'h4dee: q<=8'h03;
	15'h4def: q<=8'hd0;
	15'h4df0: q<=8'h02;
	15'h4df1: q<=8'ha9;
	15'h4df2: q<=8'h07;
	15'h4df3: q<=8'ha0;
	15'h4df4: q<=8'hff;
	15'h4df5: q<=8'hd0;
	15'h4df6: q<=8'h08;
	15'h4df7: q<=8'ha9;
	15'h4df8: q<=8'h03;
	15'h4df9: q<=8'hd0;
	15'h4dfa: q<=8'h02;
	15'h4dfb: q<=8'ha9;
	15'h4dfc: q<=8'h04;
	15'h4dfd: q<=8'ha0;
	15'h4dfe: q<=8'h00;
	15'h4dff: q<=8'h8c;
	15'h4e00: q<=8'hc6;
	15'h4e01: q<=8'h01;
	15'h4e02: q<=8'h48;
	15'h4e03: q<=8'h0d;
	15'h4e04: q<=8'hc7;
	15'h4e05: q<=8'h01;
	15'h4e06: q<=8'h8d;
	15'h4e07: q<=8'hc7;
	15'h4e08: q<=8'h01;
	15'h4e09: q<=8'h68;
	15'h4e0a: q<=8'h0d;
	15'h4e0b: q<=8'hc8;
	15'h4e0c: q<=8'h01;
	15'h4e0d: q<=8'h8d;
	15'h4e0e: q<=8'hc8;
	15'h4e0f: q<=8'h01;
	15'h4e10: q<=8'h60;
	15'h4e11: q<=8'ha9;
	15'h4e12: q<=8'h07;
	15'h4e13: q<=8'h8d;
	15'h4e14: q<=8'hc7;
	15'h4e15: q<=8'h01;
	15'h4e16: q<=8'ha9;
	15'h4e17: q<=8'h00;
	15'h4e18: q<=8'h8d;
	15'h4e19: q<=8'hc8;
	15'h4e1a: q<=8'h01;
	15'h4e1b: q<=8'had;
	15'h4e1c: q<=8'hca;
	15'h4e1d: q<=8'h01;
	15'h4e1e: q<=8'hd0;
	15'h4e1f: q<=8'h4b;
	15'h4e20: q<=8'had;
	15'h4e21: q<=8'hc7;
	15'h4e22: q<=8'h01;
	15'h4e23: q<=8'hf0;
	15'h4e24: q<=8'h46;
	15'h4e25: q<=8'ha2;
	15'h4e26: q<=8'h00;
	15'h4e27: q<=8'h8e;
	15'h4e28: q<=8'hcb;
	15'h4e29: q<=8'h01;
	15'h4e2a: q<=8'h8e;
	15'h4e2b: q<=8'hcf;
	15'h4e2c: q<=8'h01;
	15'h4e2d: q<=8'h8e;
	15'h4e2e: q<=8'hce;
	15'h4e2f: q<=8'h01;
	15'h4e30: q<=8'ha2;
	15'h4e31: q<=8'h08;
	15'h4e32: q<=8'h38;
	15'h4e33: q<=8'h6e;
	15'h4e34: q<=8'hce;
	15'h4e35: q<=8'h01;
	15'h4e36: q<=8'h0a;
	15'h4e37: q<=8'hca;
	15'h4e38: q<=8'h90;
	15'h4e39: q<=8'hf9;
	15'h4e3a: q<=8'ha0;
	15'h4e3b: q<=8'h80;
	15'h4e3c: q<=8'had;
	15'h4e3d: q<=8'hce;
	15'h4e3e: q<=8'h01;
	15'h4e3f: q<=8'h2d;
	15'h4e40: q<=8'hc8;
	15'h4e41: q<=8'h01;
	15'h4e42: q<=8'hd0;
	15'h4e43: q<=8'h02;
	15'h4e44: q<=8'ha0;
	15'h4e45: q<=8'h20;
	15'h4e46: q<=8'h8c;
	15'h4e47: q<=8'hca;
	15'h4e48: q<=8'h01;
	15'h4e49: q<=8'had;
	15'h4e4a: q<=8'hce;
	15'h4e4b: q<=8'h01;
	15'h4e4c: q<=8'h4d;
	15'h4e4d: q<=8'hc7;
	15'h4e4e: q<=8'h01;
	15'h4e4f: q<=8'h8d;
	15'h4e50: q<=8'hc7;
	15'h4e51: q<=8'h01;
	15'h4e52: q<=8'h8a;
	15'h4e53: q<=8'h0a;
	15'h4e54: q<=8'haa;
	15'h4e55: q<=8'hbd;
	15'h4e56: q<=8'hdd;
	15'h4e57: q<=8'hdd;
	15'h4e58: q<=8'h8d;
	15'h4e59: q<=8'hcc;
	15'h4e5a: q<=8'h01;
	15'h4e5b: q<=8'hbd;
	15'h4e5c: q<=8'hde;
	15'h4e5d: q<=8'hdd;
	15'h4e5e: q<=8'h8d;
	15'h4e5f: q<=8'hcd;
	15'h4e60: q<=8'h01;
	15'h4e61: q<=8'hbd;
	15'h4e62: q<=8'he3;
	15'h4e63: q<=8'hdd;
	15'h4e64: q<=8'h85;
	15'h4e65: q<=8'hbd;
	15'h4e66: q<=8'hbd;
	15'h4e67: q<=8'he4;
	15'h4e68: q<=8'hdd;
	15'h4e69: q<=8'h85;
	15'h4e6a: q<=8'hbe;
	15'h4e6b: q<=8'ha0;
	15'h4e6c: q<=8'h00;
	15'h4e6d: q<=8'h8c;
	15'h4e6e: q<=8'h40;
	15'h4e6f: q<=8'h60;
	15'h4e70: q<=8'had;
	15'h4e71: q<=8'hca;
	15'h4e72: q<=8'h01;
	15'h4e73: q<=8'hd0;
	15'h4e74: q<=8'h01;
	15'h4e75: q<=8'h60;
	15'h4e76: q<=8'hac;
	15'h4e77: q<=8'hcb;
	15'h4e78: q<=8'h01;
	15'h4e79: q<=8'hae;
	15'h4e7a: q<=8'hcc;
	15'h4e7b: q<=8'h01;
	15'h4e7c: q<=8'h0a;
	15'h4e7d: q<=8'h90;
	15'h4e7e: q<=8'h0d;
	15'h4e7f: q<=8'h9d;
	15'h4e80: q<=8'h00;
	15'h4e81: q<=8'h60;
	15'h4e82: q<=8'ha9;
	15'h4e83: q<=8'h40;
	15'h4e84: q<=8'h8d;
	15'h4e85: q<=8'hca;
	15'h4e86: q<=8'h01;
	15'h4e87: q<=8'ha0;
	15'h4e88: q<=8'h0e;
	15'h4e89: q<=8'hb8;
	15'h4e8a: q<=8'h50;
	15'h4e8b: q<=8'h73;
	15'h4e8c: q<=8'h10;
	15'h4e8d: q<=8'h25;
	15'h4e8e: q<=8'ha9;
	15'h4e8f: q<=8'h80;
	15'h4e90: q<=8'h8d;
	15'h4e91: q<=8'hca;
	15'h4e92: q<=8'h01;
	15'h4e93: q<=8'had;
	15'h4e94: q<=8'hc6;
	15'h4e95: q<=8'h01;
	15'h4e96: q<=8'hf0;
	15'h4e97: q<=8'h04;
	15'h4e98: q<=8'ha9;
	15'h4e99: q<=8'h00;
	15'h4e9a: q<=8'h91;
	15'h4e9b: q<=8'hbd;
	15'h4e9c: q<=8'hb1;
	15'h4e9d: q<=8'hbd;
	15'h4e9e: q<=8'hec;
	15'h4e9f: q<=8'hcd;
	15'h4ea0: q<=8'h01;
	15'h4ea1: q<=8'h90;
	15'h4ea2: q<=8'h08;
	15'h4ea3: q<=8'ha9;
	15'h4ea4: q<=8'h00;
	15'h4ea5: q<=8'h8d;
	15'h4ea6: q<=8'hca;
	15'h4ea7: q<=8'h01;
	15'h4ea8: q<=8'had;
	15'h4ea9: q<=8'hcf;
	15'h4eaa: q<=8'h01;
	15'h4eab: q<=8'h9d;
	15'h4eac: q<=8'h00;
	15'h4ead: q<=8'h60;
	15'h4eae: q<=8'ha0;
	15'h4eaf: q<=8'h0c;
	15'h4eb0: q<=8'hb8;
	15'h4eb1: q<=8'h50;
	15'h4eb2: q<=8'h3f;
	15'h4eb3: q<=8'ha9;
	15'h4eb4: q<=8'h08;
	15'h4eb5: q<=8'h8d;
	15'h4eb6: q<=8'h40;
	15'h4eb7: q<=8'h60;
	15'h4eb8: q<=8'h9d;
	15'h4eb9: q<=8'h00;
	15'h4eba: q<=8'h60;
	15'h4ebb: q<=8'ha9;
	15'h4ebc: q<=8'h09;
	15'h4ebd: q<=8'h8d;
	15'h4ebe: q<=8'h40;
	15'h4ebf: q<=8'h60;
	15'h4ec0: q<=8'hea;
	15'h4ec1: q<=8'ha9;
	15'h4ec2: q<=8'h08;
	15'h4ec3: q<=8'h8d;
	15'h4ec4: q<=8'h40;
	15'h4ec5: q<=8'h60;
	15'h4ec6: q<=8'hec;
	15'h4ec7: q<=8'hcd;
	15'h4ec8: q<=8'h01;
	15'h4ec9: q<=8'had;
	15'h4eca: q<=8'h50;
	15'h4ecb: q<=8'h60;
	15'h4ecc: q<=8'h90;
	15'h4ecd: q<=8'h20;
	15'h4ece: q<=8'h4d;
	15'h4ecf: q<=8'hcf;
	15'h4ed0: q<=8'h01;
	15'h4ed1: q<=8'hf0;
	15'h4ed2: q<=8'h13;
	15'h4ed3: q<=8'ha9;
	15'h4ed4: q<=8'h00;
	15'h4ed5: q<=8'hac;
	15'h4ed6: q<=8'hcb;
	15'h4ed7: q<=8'h01;
	15'h4ed8: q<=8'h91;
	15'h4ed9: q<=8'hbd;
	15'h4eda: q<=8'h88;
	15'h4edb: q<=8'h10;
	15'h4edc: q<=8'hfb;
	15'h4edd: q<=8'had;
	15'h4ede: q<=8'hce;
	15'h4edf: q<=8'h01;
	15'h4ee0: q<=8'h0d;
	15'h4ee1: q<=8'hc9;
	15'h4ee2: q<=8'h01;
	15'h4ee3: q<=8'h8d;
	15'h4ee4: q<=8'hc9;
	15'h4ee5: q<=8'h01;
	15'h4ee6: q<=8'ha9;
	15'h4ee7: q<=8'h00;
	15'h4ee8: q<=8'h8d;
	15'h4ee9: q<=8'hca;
	15'h4eea: q<=8'h01;
	15'h4eeb: q<=8'hb8;
	15'h4eec: q<=8'h50;
	15'h4eed: q<=8'h02;
	15'h4eee: q<=8'h91;
	15'h4eef: q<=8'hbd;
	15'h4ef0: q<=8'ha0;
	15'h4ef1: q<=8'h00;
	15'h4ef2: q<=8'h18;
	15'h4ef3: q<=8'h6d;
	15'h4ef4: q<=8'hcf;
	15'h4ef5: q<=8'h01;
	15'h4ef6: q<=8'h8d;
	15'h4ef7: q<=8'hcf;
	15'h4ef8: q<=8'h01;
	15'h4ef9: q<=8'hee;
	15'h4efa: q<=8'hcb;
	15'h4efb: q<=8'h01;
	15'h4efc: q<=8'hee;
	15'h4efd: q<=8'hcc;
	15'h4efe: q<=8'h01;
	15'h4eff: q<=8'h8c;
	15'h4f00: q<=8'h40;
	15'h4f01: q<=8'h60;
	15'h4f02: q<=8'h98;
	15'h4f03: q<=8'hd0;
	15'h4f04: q<=8'h03;
	15'h4f05: q<=8'h4c;
	15'h4f06: q<=8'h1b;
	15'h4f07: q<=8'hde;
	15'h4f08: q<=8'h60;
	15'h4f09: q<=8'ha9;
	15'h4f0a: q<=8'hc0;
	15'h4f0b: q<=8'hd0;
	15'h4f0c: q<=8'h05;
	15'h4f0d: q<=8'h20;
	15'h4f0e: q<=8'h53;
	15'h4f0f: q<=8'hdf;
	15'h4f10: q<=8'ha9;
	15'h4f11: q<=8'h20;
	15'h4f12: q<=8'ha0;
	15'h4f13: q<=8'h00;
	15'h4f14: q<=8'h91;
	15'h4f15: q<=8'h74;
	15'h4f16: q<=8'h4c;
	15'h4f17: q<=8'hac;
	15'h4f18: q<=8'hdf;
	15'h4f19: q<=8'h90;
	15'h4f1a: q<=8'h04;
	15'h4f1b: q<=8'h29;
	15'h4f1c: q<=8'h0f;
	15'h4f1d: q<=8'hf0;
	15'h4f1e: q<=8'h05;
	15'h4f1f: q<=8'h29;
	15'h4f20: q<=8'h0f;
	15'h4f21: q<=8'h18;
	15'h4f22: q<=8'h69;
	15'h4f23: q<=8'h01;
	15'h4f24: q<=8'h08;
	15'h4f25: q<=8'h0a;
	15'h4f26: q<=8'ha0;
	15'h4f27: q<=8'h00;
	15'h4f28: q<=8'haa;
	15'h4f29: q<=8'hbd;
	15'h4f2a: q<=8'he4;
	15'h4f2b: q<=8'h31;
	15'h4f2c: q<=8'h91;
	15'h4f2d: q<=8'h74;
	15'h4f2e: q<=8'hbd;
	15'h4f2f: q<=8'he5;
	15'h4f30: q<=8'h31;
	15'h4f31: q<=8'hc8;
	15'h4f32: q<=8'h91;
	15'h4f33: q<=8'h74;
	15'h4f34: q<=8'h20;
	15'h4f35: q<=8'h5f;
	15'h4f36: q<=8'hdf;
	15'h4f37: q<=8'h28;
	15'h4f38: q<=8'h60;
	15'h4f39: q<=8'h4a;
	15'h4f3a: q<=8'h29;
	15'h4f3b: q<=8'h0f;
	15'h4f3c: q<=8'h09;
	15'h4f3d: q<=8'ha0;
	15'h4f3e: q<=8'ha0;
	15'h4f3f: q<=8'h01;
	15'h4f40: q<=8'h91;
	15'h4f41: q<=8'h74;
	15'h4f42: q<=8'h88;
	15'h4f43: q<=8'h8a;
	15'h4f44: q<=8'h6a;
	15'h4f45: q<=8'h91;
	15'h4f46: q<=8'h74;
	15'h4f47: q<=8'hc8;
	15'h4f48: q<=8'hd0;
	15'h4f49: q<=8'h15;
	15'h4f4a: q<=8'ha4;
	15'h4f4b: q<=8'h73;
	15'h4f4c: q<=8'h09;
	15'h4f4d: q<=8'h60;
	15'h4f4e: q<=8'haa;
	15'h4f4f: q<=8'h98;
	15'h4f50: q<=8'h4c;
	15'h4f51: q<=8'h57;
	15'h4f52: q<=8'hdf;
	15'h4f53: q<=8'ha9;
	15'h4f54: q<=8'h40;
	15'h4f55: q<=8'ha2;
	15'h4f56: q<=8'h80;
	15'h4f57: q<=8'ha0;
	15'h4f58: q<=8'h00;
	15'h4f59: q<=8'h91;
	15'h4f5a: q<=8'h74;
	15'h4f5b: q<=8'hc8;
	15'h4f5c: q<=8'h8a;
	15'h4f5d: q<=8'h91;
	15'h4f5e: q<=8'h74;
	15'h4f5f: q<=8'h98;
	15'h4f60: q<=8'h38;
	15'h4f61: q<=8'h65;
	15'h4f62: q<=8'h74;
	15'h4f63: q<=8'h85;
	15'h4f64: q<=8'h74;
	15'h4f65: q<=8'h90;
	15'h4f66: q<=8'h02;
	15'h4f67: q<=8'he6;
	15'h4f68: q<=8'h75;
	15'h4f69: q<=8'h60;
	15'h4f6a: q<=8'ha0;
	15'h4f6b: q<=8'h00;
	15'h4f6c: q<=8'h09;
	15'h4f6d: q<=8'h70;
	15'h4f6e: q<=8'haa;
	15'h4f6f: q<=8'h98;
	15'h4f70: q<=8'h4c;
	15'h4f71: q<=8'h57;
	15'h4f72: q<=8'hdf;
	15'h4f73: q<=8'h84;
	15'h4f74: q<=8'h73;
	15'h4f75: q<=8'ha0;
	15'h4f76: q<=8'h00;
	15'h4f77: q<=8'h0a;
	15'h4f78: q<=8'h90;
	15'h4f79: q<=8'h01;
	15'h4f7a: q<=8'h88;
	15'h4f7b: q<=8'h84;
	15'h4f7c: q<=8'h6f;
	15'h4f7d: q<=8'h0a;
	15'h4f7e: q<=8'h26;
	15'h4f7f: q<=8'h6f;
	15'h4f80: q<=8'h85;
	15'h4f81: q<=8'h6e;
	15'h4f82: q<=8'h8a;
	15'h4f83: q<=8'h0a;
	15'h4f84: q<=8'ha0;
	15'h4f85: q<=8'h00;
	15'h4f86: q<=8'h90;
	15'h4f87: q<=8'h01;
	15'h4f88: q<=8'h88;
	15'h4f89: q<=8'h84;
	15'h4f8a: q<=8'h71;
	15'h4f8b: q<=8'h0a;
	15'h4f8c: q<=8'h26;
	15'h4f8d: q<=8'h71;
	15'h4f8e: q<=8'h85;
	15'h4f8f: q<=8'h70;
	15'h4f90: q<=8'ha2;
	15'h4f91: q<=8'h6e;
	15'h4f92: q<=8'ha0;
	15'h4f93: q<=8'h00;
	15'h4f94: q<=8'hb5;
	15'h4f95: q<=8'h02;
	15'h4f96: q<=8'h91;
	15'h4f97: q<=8'h74;
	15'h4f98: q<=8'hb5;
	15'h4f99: q<=8'h03;
	15'h4f9a: q<=8'h29;
	15'h4f9b: q<=8'h1f;
	15'h4f9c: q<=8'hc8;
	15'h4f9d: q<=8'h91;
	15'h4f9e: q<=8'h74;
	15'h4f9f: q<=8'hb5;
	15'h4fa0: q<=8'h00;
	15'h4fa1: q<=8'hc8;
	15'h4fa2: q<=8'h91;
	15'h4fa3: q<=8'h74;
	15'h4fa4: q<=8'hb5;
	15'h4fa5: q<=8'h01;
	15'h4fa6: q<=8'h45;
	15'h4fa7: q<=8'h73;
	15'h4fa8: q<=8'h29;
	15'h4fa9: q<=8'h1f;
	15'h4faa: q<=8'h45;
	15'h4fab: q<=8'h73;
	15'h4fac: q<=8'hc8;
	15'h4fad: q<=8'h91;
	15'h4fae: q<=8'h74;
	15'h4faf: q<=8'hd0;
	15'h4fb0: q<=8'hae;
	15'h4fb1: q<=8'h38;
	15'h4fb2: q<=8'h08;
	15'h4fb3: q<=8'h88;
	15'h4fb4: q<=8'h84;
	15'h4fb5: q<=8'hae;
	15'h4fb6: q<=8'h18;
	15'h4fb7: q<=8'h65;
	15'h4fb8: q<=8'hae;
	15'h4fb9: q<=8'h28;
	15'h4fba: q<=8'haa;
	15'h4fbb: q<=8'h08;
	15'h4fbc: q<=8'h86;
	15'h4fbd: q<=8'haf;
	15'h4fbe: q<=8'hb5;
	15'h4fbf: q<=8'h00;
	15'h4fc0: q<=8'h4a;
	15'h4fc1: q<=8'h4a;
	15'h4fc2: q<=8'h4a;
	15'h4fc3: q<=8'h4a;
	15'h4fc4: q<=8'h28;
	15'h4fc5: q<=8'h20;
	15'h4fc6: q<=8'h19;
	15'h4fc7: q<=8'hdf;
	15'h4fc8: q<=8'ha5;
	15'h4fc9: q<=8'hae;
	15'h4fca: q<=8'hd0;
	15'h4fcb: q<=8'h01;
	15'h4fcc: q<=8'h18;
	15'h4fcd: q<=8'ha6;
	15'h4fce: q<=8'haf;
	15'h4fcf: q<=8'hb5;
	15'h4fd0: q<=8'h00;
	15'h4fd1: q<=8'h20;
	15'h4fd2: q<=8'h19;
	15'h4fd3: q<=8'hdf;
	15'h4fd4: q<=8'ha6;
	15'h4fd5: q<=8'haf;
	15'h4fd6: q<=8'hca;
	15'h4fd7: q<=8'hc6;
	15'h4fd8: q<=8'hae;
	15'h4fd9: q<=8'h10;
	15'h4fda: q<=8'he0;
	15'h4fdb: q<=8'h60;
	15'h4fdc: q<=8'h10;
	15'h4fdd: q<=8'h10;
	15'h4fde: q<=8'h40;
	15'h4fdf: q<=8'h40;
	15'h4fe0: q<=8'h90;
	15'h4fe1: q<=8'h90;
	15'h4fe2: q<=8'hff;
	15'h4fe3: q<=8'hff;
	15'h4fe4: q<=8'h00;
	15'h4fe5: q<=8'h0c;
	15'h4fe6: q<=8'h16;
	15'h4fe7: q<=8'h1e;
	15'h4fe8: q<=8'h20;
	15'h4fe9: q<=8'h1e;
	15'h4fea: q<=8'h16;
	15'h4feb: q<=8'h0c;
	15'h4fec: q<=8'h00;
	15'h4fed: q<=8'hf4;
	15'h4fee: q<=8'hea;
	15'h4fef: q<=8'he2;
	15'h4ff0: q<=8'he0;
	15'h4ff1: q<=8'he2;
	15'h4ff2: q<=8'hea;
	15'h4ff3: q<=8'hf4;
	15'h4ff4: q<=8'h00;
	15'h4ff5: q<=8'h0c;
	15'h4ff6: q<=8'h16;
	15'h4ff7: q<=8'h1e;
	15'h4ff8: q<=8'h00;
	15'h4ff9: q<=8'h00;
	15'h4ffa: q<=8'h04;
	15'h4ffb: q<=8'hd7;
	15'h4ffc: q<=8'h3f;
	15'h4ffd: q<=8'hd9;
	15'h4ffe: q<=8'h04;
	15'h4fff: q<=8'hd7;
	15'h5000: q<=8'he6;
	15'h5001: q<=8'h06;
	15'h5002: q<=8'h85;
	15'h5003: q<=8'h17;
	15'h5004: q<=8'ha5;
	15'h5005: q<=8'h07;
	15'h5006: q<=8'h4a;
	15'h5007: q<=8'hb0;
	15'h5008: q<=8'h27;
	15'h5009: q<=8'ha0;
	15'h500a: q<=8'h00;
	15'h500b: q<=8'ha2;
	15'h500c: q<=8'h02;
	15'h500d: q<=8'hb5;
	15'h500e: q<=8'h13;
	15'h500f: q<=8'hf0;
	15'h5010: q<=8'h09;
	15'h5011: q<=8'hc9;
	15'h5012: q<=8'h10;
	15'h5013: q<=8'h90;
	15'h5014: q<=8'h05;
	15'h5015: q<=8'h69;
	15'h5016: q<=8'hef;
	15'h5017: q<=8'hc8;
	15'h5018: q<=8'h95;
	15'h5019: q<=8'h13;
	15'h501a: q<=8'hca;
	15'h501b: q<=8'h10;
	15'h501c: q<=8'hf0;
	15'h501d: q<=8'h98;
	15'h501e: q<=8'hd0;
	15'h501f: q<=8'h10;
	15'h5020: q<=8'ha2;
	15'h5021: q<=8'h02;
	15'h5022: q<=8'hb5;
	15'h5023: q<=8'h13;
	15'h5024: q<=8'hf0;
	15'h5025: q<=8'h07;
	15'h5026: q<=8'h18;
	15'h5027: q<=8'h69;
	15'h5028: q<=8'hef;
	15'h5029: q<=8'h95;
	15'h502a: q<=8'h13;
	15'h502b: q<=8'h30;
	15'h502c: q<=8'h03;
	15'h502d: q<=8'hca;
	15'h502e: q<=8'h10;
	15'h502f: q<=8'hf2;
	15'h5030: q<=8'h60;
	15'h5031: q<=8'h5d;
	15'h5032: q<=8'hd1;
	15'h5033: q<=8'h8f;
	15'h5034: q<=8'hd1;
	15'h5035: q<=8'h8f;
	15'h5036: q<=8'hd1;
	15'h5037: q<=8'hb1;
	15'h5038: q<=8'hd1;
	15'h5039: q<=8'heb;
	15'h503a: q<=8'hd1;
	15'h503b: q<=8'h03;
	15'h503c: q<=8'hd2;
	15'h503d: q<=8'h61;
	15'h503e: q<=8'hd2;
	15'h503f: q<=8'hcb;
	15'h5040: q<=8'hd2;
	15'h5041: q<=8'h33;
	15'h5042: q<=8'hd3;
	15'h5043: q<=8'h66;
	15'h5044: q<=8'hd3;
	15'h5045: q<=8'hb0;
	15'h5046: q<=8'hd3;
	15'h5047: q<=8'he6;
	15'h5048: q<=8'hd3;
	15'h5049: q<=8'hff;
	15'h504a: q<=8'hd3;
	15'h504b: q<=8'h17;
	15'h504c: q<=8'hd4;
	15'h504d: q<=8'h1d;
	15'h504e: q<=8'hd4;
	15'h504f: q<=8'h34;
	15'h5050: q<=8'hd4;
	15'h5051: q<=8'h4c;
	15'h5052: q<=8'hd4;
	15'h5053: q<=8'h60;
	15'h5054: q<=8'hd4;
	15'h5055: q<=8'ha1;
	15'h5056: q<=8'hd4;
	15'h5057: q<=8'hab;
	15'h5058: q<=8'hd4;
	15'h5059: q<=8'hef;
	15'h505a: q<=8'hd4;
	15'h505b: q<=8'h30;
	15'h505c: q<=8'hd5;
	15'h505d: q<=8'h75;
	15'h505e: q<=8'hd5;
	15'h505f: q<=8'h85;
	15'h5060: q<=8'hd5;
	15'h5061: q<=8'ha1;
	15'h5062: q<=8'hd5;
	15'h5063: q<=8'ha8;
	15'h5064: q<=8'hd5;
	15'h5065: q<=8'he9;
	15'h5066: q<=8'hd5;
	15'h5067: q<=8'h1c;
	15'h5068: q<=8'hd6;
	15'h5069: q<=8'h62;
	15'h506a: q<=8'hd6;
	15'h506b: q<=8'h7a;
	15'h506c: q<=8'hd6;
	15'h506d: q<=8'h67;
	15'h506e: q<=8'hd1;
	15'h506f: q<=8'h97;
	15'h5070: q<=8'hd1;
	15'h5071: q<=8'h97;
	15'h5072: q<=8'hd1;
	15'h5073: q<=8'hbd;
	15'h5074: q<=8'hd1;
	15'h5075: q<=8'hf0;
	15'h5076: q<=8'hd1;
	15'h5077: q<=8'h17;
	15'h5078: q<=8'hd2;
	15'h5079: q<=8'h75;
	15'h507a: q<=8'hd2;
	15'h507b: q<=8'he0;
	15'h507c: q<=8'hd2;
	15'h507d: q<=8'h3f;
	15'h507e: q<=8'hd3;
	15'h507f: q<=8'h79;
	15'h5080: q<=8'hd3;
	15'h5081: q<=8'hbe;
	15'h5082: q<=8'hd3;
	15'h5083: q<=8'he6;
	15'h5084: q<=8'hd3;
	15'h5085: q<=8'hff;
	15'h5086: q<=8'hd3;
	15'h5087: q<=8'h17;
	15'h5088: q<=8'hd4;
	15'h5089: q<=8'h22;
	15'h508a: q<=8'hd4;
	15'h508b: q<=8'h3a;
	15'h508c: q<=8'hd4;
	15'h508d: q<=8'h51;
	15'h508e: q<=8'hd4;
	15'h508f: q<=8'h6d;
	15'h5090: q<=8'hd4;
	15'h5091: q<=8'ha1;
	15'h5092: q<=8'hd4;
	15'h5093: q<=8'hba;
	15'h5094: q<=8'hd4;
	15'h5095: q<=8'hfd;
	15'h5096: q<=8'hd4;
	15'h5097: q<=8'h3f;
	15'h5098: q<=8'hd5;
	15'h5099: q<=8'h75;
	15'h509a: q<=8'hd5;
	15'h509b: q<=8'h85;
	15'h509c: q<=8'hd5;
	15'h509d: q<=8'ha1;
	15'h509e: q<=8'hd5;
	15'h509f: q<=8'hb9;
	15'h50a0: q<=8'hd5;
	15'h50a1: q<=8'hf6;
	15'h50a2: q<=8'hd5;
	15'h50a3: q<=8'h29;
	15'h50a4: q<=8'hd6;
	15'h50a5: q<=8'h68;
	15'h50a6: q<=8'hd6;
	15'h50a7: q<=8'h7a;
	15'h50a8: q<=8'hd6;
	15'h50a9: q<=8'h75;
	15'h50aa: q<=8'hd1;
	15'h50ab: q<=8'h9f;
	15'h50ac: q<=8'hd1;
	15'h50ad: q<=8'h9f;
	15'h50ae: q<=8'hd1;
	15'h50af: q<=8'hcf;
	15'h50b0: q<=8'hd1;
	15'h50b1: q<=8'hf6;
	15'h50b2: q<=8'hd1;
	15'h50b3: q<=8'h30;
	15'h50b4: q<=8'hd2;
	15'h50b5: q<=8'h94;
	15'h50b6: q<=8'hd2;
	15'h50b7: q<=8'hfb;
	15'h50b8: q<=8'hd2;
	15'h50b9: q<=8'h50;
	15'h50ba: q<=8'hd3;
	15'h50bb: q<=8'h8b;
	15'h50bc: q<=8'hd3;
	15'h50bd: q<=8'hcb;
	15'h50be: q<=8'hd3;
	15'h50bf: q<=8'hf5;
	15'h50c0: q<=8'hd3;
	15'h50c1: q<=8'h0e;
	15'h50c2: q<=8'hd4;
	15'h50c3: q<=8'h17;
	15'h50c4: q<=8'hd4;
	15'h50c5: q<=8'h28;
	15'h50c6: q<=8'hd4;
	15'h50c7: q<=8'h41;
	15'h50c8: q<=8'hd4;
	15'h50c9: q<=8'h5b;
	15'h50ca: q<=8'hd4;
	15'h50cb: q<=8'h83;
	15'h50cc: q<=8'hd4;
	15'h50cd: q<=8'ha1;
	15'h50ce: q<=8'hd4;
	15'h50cf: q<=8'hcc;
	15'h50d0: q<=8'hd4;
	15'h50d1: q<=8'h0e;
	15'h50d2: q<=8'hd5;
	15'h50d3: q<=8'h51;
	15'h50d4: q<=8'hd5;
	15'h50d5: q<=8'h75;
	15'h50d6: q<=8'hd5;
	15'h50d7: q<=8'h8e;
	15'h50d8: q<=8'hd5;
	15'h50d9: q<=8'ha1;
	15'h50da: q<=8'hd5;
	15'h50db: q<=8'hc8;
	15'h50dc: q<=8'hd5;
	15'h50dd: q<=8'h04;
	15'h50de: q<=8'hd6;
	15'h50df: q<=8'h3e;
	15'h50e0: q<=8'hd6;
	15'h50e1: q<=8'h6f;
	15'h50e2: q<=8'hd6;
	15'h50e3: q<=8'h8f;
	15'h50e4: q<=8'hd6;
	15'h50e5: q<=8'h7f;
	15'h50e6: q<=8'hd1;
	15'h50e7: q<=8'ha8;
	15'h50e8: q<=8'hd1;
	15'h50e9: q<=8'ha8;
	15'h50ea: q<=8'hd1;
	15'h50eb: q<=8'hde;
	15'h50ec: q<=8'hd1;
	15'h50ed: q<=8'hfc;
	15'h50ee: q<=8'hd1;
	15'h50ef: q<=8'h4d;
	15'h50f0: q<=8'hd2;
	15'h50f1: q<=8'hae;
	15'h50f2: q<=8'hd2;
	15'h50f3: q<=8'h16;
	15'h50f4: q<=8'hd3;
	15'h50f5: q<=8'h5e;
	15'h50f6: q<=8'hd3;
	15'h50f7: q<=8'ha0;
	15'h50f8: q<=8'hd3;
	15'h50f9: q<=8'hda;
	15'h50fa: q<=8'hd3;
	15'h50fb: q<=8'hed;
	15'h50fc: q<=8'hd3;
	15'h50fd: q<=8'h06;
	15'h50fe: q<=8'hd4;
	15'h50ff: q<=8'h17;
	15'h5100: q<=8'hd4;
	15'h5101: q<=8'h2d;
	15'h5102: q<=8'hd4;
	15'h5103: q<=8'h46;
	15'h5104: q<=8'hd4;
	15'h5105: q<=8'h56;
	15'h5106: q<=8'hd4;
	15'h5107: q<=8'h92;
	15'h5108: q<=8'hd4;
	15'h5109: q<=8'ha1;
	15'h510a: q<=8'hd4;
	15'h510b: q<=8'hdd;
	15'h510c: q<=8'hd4;
	15'h510d: q<=8'h1f;
	15'h510e: q<=8'hd5;
	15'h510f: q<=8'h63;
	15'h5110: q<=8'hd5;
	15'h5111: q<=8'h75;
	15'h5112: q<=8'hd5;
	15'h5113: q<=8'h97;
	15'h5114: q<=8'hd5;
	15'h5115: q<=8'ha1;
	15'h5116: q<=8'hd5;
	15'h5117: q<=8'hd9;
	15'h5118: q<=8'hd5;
	15'h5119: q<=8'h10;
	15'h511a: q<=8'hd6;
	15'h511b: q<=8'h51;
	15'h511c: q<=8'hd6;
	15'h511d: q<=8'h74;
	15'h511e: q<=8'hd6;
	15'h511f: q<=8'ha1;
	15'h5120: q<=8'hd6;
	15'h5121: q<=8'h51;
	15'h5122: q<=8'h56;
	15'h5123: q<=8'h00;
	15'h5124: q<=8'h1a;
	15'h5125: q<=8'h01;
	15'h5126: q<=8'h20;
	15'h5127: q<=8'h31;
	15'h5128: q<=8'h56;
	15'h5129: q<=8'h01;
	15'h512a: q<=8'h38;
	15'h512b: q<=8'h31;
	15'h512c: q<=8'hb0;
	15'h512d: q<=8'h41;
	15'h512e: q<=8'h00;
	15'h512f: q<=8'h11;
	15'h5130: q<=8'hf6;
	15'h5131: q<=8'h30;
	15'h5132: q<=8'h38;
	15'h5133: q<=8'h31;
	15'h5134: q<=8'hce;
	15'h5135: q<=8'h51;
	15'h5136: q<=8'h0a;
	15'h5137: q<=8'h31;
	15'h5138: q<=8'he2;
	15'h5139: q<=8'h31;
	15'h513a: q<=8'he2;
	15'h513b: q<=8'h51;
	15'h513c: q<=8'hba;
	15'h513d: q<=8'h51;
	15'h513e: q<=8'h98;
	15'h513f: q<=8'h51;
	15'h5140: q<=8'hd8;
	15'h5141: q<=8'h51;
	15'h5142: q<=8'hc9;
	15'h5143: q<=8'h31;
	15'h5144: q<=8'h56;
	15'h5145: q<=8'h51;
	15'h5146: q<=8'h80;
	15'h5147: q<=8'h51;
	15'h5148: q<=8'h80;
	15'h5149: q<=8'h51;
	15'h514a: q<=8'h80;
	15'h514b: q<=8'h51;
	15'h514c: q<=8'h80;
	15'h514d: q<=8'h71;
	15'h514e: q<=8'h92;
	15'h514f: q<=8'h51;
	15'h5150: q<=8'h80;
	15'h5151: q<=8'h31;
	15'h5152: q<=8'hb0;
	15'h5153: q<=8'h51;
	15'h5154: q<=8'h89;
	15'h5155: q<=8'h41;
	15'h5156: q<=8'h89;
	15'h5157: q<=8'h00;
	15'h5158: q<=8'h00;
	15'h5159: q<=8'h71;
	15'h515a: q<=8'h5a;
	15'h515b: q<=8'h71;
	15'h515c: q<=8'ha0;
	15'h515d: q<=8'he5;
	15'h515e: q<=8'h22;
	15'h515f: q<=8'h16;
	15'h5160: q<=8'h2e;
	15'h5161: q<=8'h1e;
	15'h5162: q<=8'h00;
	15'h5163: q<=8'h32;
	15'h5164: q<=8'h40;
	15'h5165: q<=8'h1e;
	15'h5166: q<=8'hb8;
	15'h5167: q<=8'hd9;
	15'h5168: q<=8'h20;
	15'h5169: q<=8'h26;
	15'h516a: q<=8'h30;
	15'h516b: q<=8'h00;
	15'h516c: q<=8'h1c;
	15'h516d: q<=8'h1e;
	15'h516e: q<=8'h00;
	15'h516f: q<=8'h34;
	15'h5170: q<=8'h16;
	15'h5171: q<=8'h38;
	15'h5172: q<=8'h3c;
	15'h5173: q<=8'h26;
	15'h5174: q<=8'h9e;
	15'h5175: q<=8'he5;
	15'h5176: q<=8'h3a;
	15'h5177: q<=8'h34;
	15'h5178: q<=8'h26;
	15'h5179: q<=8'h1e;
	15'h517a: q<=8'h2c;
	15'h517b: q<=8'h1e;
	15'h517c: q<=8'h30;
	15'h517d: q<=8'h1c;
	15'h517e: q<=8'h9e;
	15'h517f: q<=8'hd3;
	15'h5180: q<=8'h28;
	15'h5181: q<=8'h3e;
	15'h5182: q<=8'h1e;
	15'h5183: q<=8'h22;
	15'h5184: q<=8'h32;
	15'h5185: q<=8'h00;
	15'h5186: q<=8'h3c;
	15'h5187: q<=8'h1e;
	15'h5188: q<=8'h38;
	15'h5189: q<=8'h2e;
	15'h518a: q<=8'h26;
	15'h518b: q<=8'h30;
	15'h518c: q<=8'h16;
	15'h518d: q<=8'h1c;
	15'h518e: q<=8'hb2;
	15'h518f: q<=8'hcd;
	15'h5190: q<=8'h34;
	15'h5191: q<=8'h2c;
	15'h5192: q<=8'h16;
	15'h5193: q<=8'h46;
	15'h5194: q<=8'h1e;
	15'h5195: q<=8'h38;
	15'h5196: q<=8'h80;
	15'h5197: q<=8'hc6;
	15'h5198: q<=8'h28;
	15'h5199: q<=8'h32;
	15'h519a: q<=8'h3e;
	15'h519b: q<=8'h1e;
	15'h519c: q<=8'h3e;
	15'h519d: q<=8'h38;
	15'h519e: q<=8'h80;
	15'h519f: q<=8'hc6;
	15'h51a0: q<=8'h3a;
	15'h51a1: q<=8'h34;
	15'h51a2: q<=8'h26;
	15'h51a3: q<=8'h1e;
	15'h51a4: q<=8'h2c;
	15'h51a5: q<=8'h1e;
	15'h51a6: q<=8'h38;
	15'h51a7: q<=8'h80;
	15'h51a8: q<=8'hc6;
	15'h51a9: q<=8'h28;
	15'h51aa: q<=8'h3e;
	15'h51ab: q<=8'h22;
	15'h51ac: q<=8'h16;
	15'h51ad: q<=8'h1c;
	15'h51ae: q<=8'h32;
	15'h51af: q<=8'h38;
	15'h51b0: q<=8'h80;
	15'h51b1: q<=8'hdf;
	15'h51b2: q<=8'h34;
	15'h51b3: q<=8'h38;
	15'h51b4: q<=8'h1e;
	15'h51b5: q<=8'h3a;
	15'h51b6: q<=8'h3a;
	15'h51b7: q<=8'h00;
	15'h51b8: q<=8'h3a;
	15'h51b9: q<=8'h3c;
	15'h51ba: q<=8'h16;
	15'h51bb: q<=8'h38;
	15'h51bc: q<=8'hbc;
	15'h51bd: q<=8'hcd;
	15'h51be: q<=8'h16;
	15'h51bf: q<=8'h34;
	15'h51c0: q<=8'h34;
	15'h51c1: q<=8'h3e;
	15'h51c2: q<=8'h46;
	15'h51c3: q<=8'h1e;
	15'h51c4: q<=8'h48;
	15'h51c5: q<=8'h00;
	15'h51c6: q<=8'h3a;
	15'h51c7: q<=8'h3e;
	15'h51c8: q<=8'h38;
	15'h51c9: q<=8'h00;
	15'h51ca: q<=8'h3a;
	15'h51cb: q<=8'h3c;
	15'h51cc: q<=8'h16;
	15'h51cd: q<=8'h38;
	15'h51ce: q<=8'hbc;
	15'h51cf: q<=8'hd6;
	15'h51d0: q<=8'h3a;
	15'h51d1: q<=8'h3c;
	15'h51d2: q<=8'h16;
	15'h51d3: q<=8'h38;
	15'h51d4: q<=8'h3c;
	15'h51d5: q<=8'h00;
	15'h51d6: q<=8'h1c;
	15'h51d7: q<=8'h38;
	15'h51d8: q<=8'h3e;
	15'h51d9: q<=8'h1e;
	15'h51da: q<=8'h1a;
	15'h51db: q<=8'h2a;
	15'h51dc: q<=8'h1e;
	15'h51dd: q<=8'hb0;
	15'h51de: q<=8'hdc;
	15'h51df: q<=8'h34;
	15'h51e0: q<=8'h3e;
	15'h51e1: q<=8'h2c;
	15'h51e2: q<=8'h3a;
	15'h51e3: q<=8'h16;
	15'h51e4: q<=8'h38;
	15'h51e5: q<=8'h00;
	15'h51e6: q<=8'h3a;
	15'h51e7: q<=8'h3c;
	15'h51e8: q<=8'h16;
	15'h51e9: q<=8'h38;
	15'h51ea: q<=8'hbc;
	15'h51eb: q<=8'hf4;
	15'h51ec: q<=8'h34;
	15'h51ed: q<=8'h2c;
	15'h51ee: q<=8'h16;
	15'h51ef: q<=8'hc6;
	15'h51f0: q<=8'hf1;
	15'h51f1: q<=8'h28;
	15'h51f2: q<=8'h32;
	15'h51f3: q<=8'h3e;
	15'h51f4: q<=8'h1e;
	15'h51f5: q<=8'hc8;
	15'h51f6: q<=8'hf1;
	15'h51f7: q<=8'h3a;
	15'h51f8: q<=8'h34;
	15'h51f9: q<=8'h26;
	15'h51fa: q<=8'h1e;
	15'h51fb: q<=8'hac;
	15'h51fc: q<=8'hee;
	15'h51fd: q<=8'h28;
	15'h51fe: q<=8'h3e;
	15'h51ff: q<=8'h1e;
	15'h5200: q<=8'h22;
	15'h5201: q<=8'h3e;
	15'h5202: q<=8'h9e;
	15'h5203: q<=8'hc7;
	15'h5204: q<=8'h1e;
	15'h5205: q<=8'h30;
	15'h5206: q<=8'h3c;
	15'h5207: q<=8'h1e;
	15'h5208: q<=8'h38;
	15'h5209: q<=8'h00;
	15'h520a: q<=8'h46;
	15'h520b: q<=8'h32;
	15'h520c: q<=8'h3e;
	15'h520d: q<=8'h38;
	15'h520e: q<=8'h00;
	15'h520f: q<=8'h26;
	15'h5210: q<=8'h30;
	15'h5211: q<=8'h26;
	15'h5212: q<=8'h3c;
	15'h5213: q<=8'h26;
	15'h5214: q<=8'h16;
	15'h5215: q<=8'h2c;
	15'h5216: q<=8'hba;
	15'h5217: q<=8'hb8;
	15'h5218: q<=8'h3a;
	15'h5219: q<=8'h40;
	15'h521a: q<=8'h34;
	15'h521b: q<=8'h00;
	15'h521c: q<=8'h1e;
	15'h521d: q<=8'h30;
	15'h521e: q<=8'h3c;
	15'h521f: q<=8'h38;
	15'h5220: q<=8'h1e;
	15'h5221: q<=8'h48;
	15'h5222: q<=8'h00;
	15'h5223: q<=8'h40;
	15'h5224: q<=8'h32;
	15'h5225: q<=8'h3a;
	15'h5226: q<=8'h00;
	15'h5227: q<=8'h26;
	15'h5228: q<=8'h30;
	15'h5229: q<=8'h26;
	15'h522a: q<=8'h3c;
	15'h522b: q<=8'h26;
	15'h522c: q<=8'h16;
	15'h522d: q<=8'h2c;
	15'h522e: q<=8'h1e;
	15'h522f: q<=8'hba;
	15'h5230: q<=8'hac;
	15'h5231: q<=8'h22;
	15'h5232: q<=8'h1e;
	15'h5233: q<=8'h18;
	15'h5234: q<=8'h1e;
	15'h5235: q<=8'h30;
	15'h5236: q<=8'h00;
	15'h5237: q<=8'h3a;
	15'h5238: q<=8'h26;
	15'h5239: q<=8'h1e;
	15'h523a: q<=8'h00;
	15'h523b: q<=8'h26;
	15'h523c: q<=8'h24;
	15'h523d: q<=8'h38;
	15'h523e: q<=8'h1e;
	15'h523f: q<=8'h00;
	15'h5240: q<=8'h26;
	15'h5241: q<=8'h30;
	15'h5242: q<=8'h26;
	15'h5243: q<=8'h3c;
	15'h5244: q<=8'h26;
	15'h5245: q<=8'h16;
	15'h5246: q<=8'h2c;
	15'h5247: q<=8'h1e;
	15'h5248: q<=8'h30;
	15'h5249: q<=8'h00;
	15'h524a: q<=8'h1e;
	15'h524b: q<=8'h26;
	15'h524c: q<=8'hb0;
	15'h524d: q<=8'hc7;
	15'h524e: q<=8'h1e;
	15'h524f: q<=8'h30;
	15'h5250: q<=8'h3c;
	15'h5251: q<=8'h38;
	15'h5252: q<=8'h1e;
	15'h5253: q<=8'h00;
	15'h5254: q<=8'h3a;
	15'h5255: q<=8'h3e;
	15'h5256: q<=8'h3a;
	15'h5257: q<=8'h00;
	15'h5258: q<=8'h26;
	15'h5259: q<=8'h30;
	15'h525a: q<=8'h26;
	15'h525b: q<=8'h1a;
	15'h525c: q<=8'h26;
	15'h525d: q<=8'h16;
	15'h525e: q<=8'h2c;
	15'h525f: q<=8'h1e;
	15'h5260: q<=8'hba;
	15'h5261: q<=8'hc7;
	15'h5262: q<=8'h3a;
	15'h5263: q<=8'h34;
	15'h5264: q<=8'h26;
	15'h5265: q<=8'h30;
	15'h5266: q<=8'h00;
	15'h5267: q<=8'h2a;
	15'h5268: q<=8'h30;
	15'h5269: q<=8'h32;
	15'h526a: q<=8'h18;
	15'h526b: q<=8'h00;
	15'h526c: q<=8'h3c;
	15'h526d: q<=8'h32;
	15'h526e: q<=8'h00;
	15'h526f: q<=8'h1a;
	15'h5270: q<=8'h24;
	15'h5271: q<=8'h16;
	15'h5272: q<=8'h30;
	15'h5273: q<=8'h22;
	15'h5274: q<=8'h9e;
	15'h5275: q<=8'ha6;
	15'h5276: q<=8'h3c;
	15'h5277: q<=8'h32;
	15'h5278: q<=8'h3e;
	15'h5279: q<=8'h38;
	15'h527a: q<=8'h30;
	15'h527b: q<=8'h1e;
	15'h527c: q<=8'h48;
	15'h527d: q<=8'h00;
	15'h527e: q<=8'h2c;
	15'h527f: q<=8'h1e;
	15'h5280: q<=8'h00;
	15'h5281: q<=8'h18;
	15'h5282: q<=8'h32;
	15'h5283: q<=8'h3e;
	15'h5284: q<=8'h3c;
	15'h5285: q<=8'h32;
	15'h5286: q<=8'h30;
	15'h5287: q<=8'h00;
	15'h5288: q<=8'h34;
	15'h5289: q<=8'h32;
	15'h528a: q<=8'h3e;
	15'h528b: q<=8'h38;
	15'h528c: q<=8'h00;
	15'h528d: q<=8'h1a;
	15'h528e: q<=8'h24;
	15'h528f: q<=8'h16;
	15'h5290: q<=8'h30;
	15'h5291: q<=8'h22;
	15'h5292: q<=8'h1e;
	15'h5293: q<=8'hb8;
	15'h5294: q<=8'hb5;
	15'h5295: q<=8'h2a;
	15'h5296: q<=8'h30;
	15'h5297: q<=8'h32;
	15'h5298: q<=8'h34;
	15'h5299: q<=8'h20;
	15'h529a: q<=8'h00;
	15'h529b: q<=8'h1c;
	15'h529c: q<=8'h38;
	15'h529d: q<=8'h1e;
	15'h529e: q<=8'h24;
	15'h529f: q<=8'h1e;
	15'h52a0: q<=8'h30;
	15'h52a1: q<=8'h00;
	15'h52a2: q<=8'h48;
	15'h52a3: q<=8'h3e;
	15'h52a4: q<=8'h2e;
	15'h52a5: q<=8'h00;
	15'h52a6: q<=8'h42;
	15'h52a7: q<=8'h1e;
	15'h52a8: q<=8'h1a;
	15'h52a9: q<=8'h24;
	15'h52aa: q<=8'h3a;
	15'h52ab: q<=8'h1e;
	15'h52ac: q<=8'h2c;
	15'h52ad: q<=8'hb0;
	15'h52ae: q<=8'hac;
	15'h52af: q<=8'h22;
	15'h52b0: q<=8'h26;
	15'h52b1: q<=8'h38;
	15'h52b2: q<=8'h1e;
	15'h52b3: q<=8'h00;
	15'h52b4: q<=8'h2c;
	15'h52b5: q<=8'h16;
	15'h52b6: q<=8'h00;
	15'h52b7: q<=8'h34;
	15'h52b8: q<=8'h1e;
	15'h52b9: q<=8'h38;
	15'h52ba: q<=8'h26;
	15'h52bb: q<=8'h2c;
	15'h52bc: q<=8'h2c;
	15'h52bd: q<=8'h16;
	15'h52be: q<=8'h00;
	15'h52bf: q<=8'h34;
	15'h52c0: q<=8'h16;
	15'h52c1: q<=8'h38;
	15'h52c2: q<=8'h16;
	15'h52c3: q<=8'h00;
	15'h52c4: q<=8'h1a;
	15'h52c5: q<=8'h16;
	15'h52c6: q<=8'h2e;
	15'h52c7: q<=8'h18;
	15'h52c8: q<=8'h26;
	15'h52c9: q<=8'h16;
	15'h52ca: q<=8'hb8;
	15'h52cb: q<=8'hc4;
	15'h52cc: q<=8'h34;
	15'h52cd: q<=8'h38;
	15'h52ce: q<=8'h1e;
	15'h52cf: q<=8'h3a;
	15'h52d0: q<=8'h3a;
	15'h52d1: q<=8'h00;
	15'h52d2: q<=8'h20;
	15'h52d3: q<=8'h26;
	15'h52d4: q<=8'h38;
	15'h52d5: q<=8'h1e;
	15'h52d6: q<=8'h00;
	15'h52d7: q<=8'h3c;
	15'h52d8: q<=8'h32;
	15'h52d9: q<=8'h00;
	15'h52da: q<=8'h3a;
	15'h52db: q<=8'h1e;
	15'h52dc: q<=8'h2c;
	15'h52dd: q<=8'h1e;
	15'h52de: q<=8'h1a;
	15'h52df: q<=8'hbc;
	15'h52e0: q<=8'hb2;
	15'h52e1: q<=8'h34;
	15'h52e2: q<=8'h32;
	15'h52e3: q<=8'h3e;
	15'h52e4: q<=8'h3a;
	15'h52e5: q<=8'h3a;
	15'h52e6: q<=8'h1e;
	15'h52e7: q<=8'h48;
	15'h52e8: q<=8'h00;
	15'h52e9: q<=8'h20;
	15'h52ea: q<=8'h1e;
	15'h52eb: q<=8'h3e;
	15'h52ec: q<=8'h00;
	15'h52ed: q<=8'h36;
	15'h52ee: q<=8'h3e;
	15'h52ef: q<=8'h16;
	15'h52f0: q<=8'h30;
	15'h52f1: q<=8'h1c;
	15'h52f2: q<=8'h00;
	15'h52f3: q<=8'h1a;
	15'h52f4: q<=8'h32;
	15'h52f5: q<=8'h38;
	15'h52f6: q<=8'h38;
	15'h52f7: q<=8'h1e;
	15'h52f8: q<=8'h1a;
	15'h52f9: q<=8'h3c;
	15'h52fa: q<=8'h9e;
	15'h52fb: q<=8'hb2;
	15'h52fc: q<=8'h20;
	15'h52fd: q<=8'h26;
	15'h52fe: q<=8'h38;
	15'h52ff: q<=8'h1e;
	15'h5300: q<=8'h00;
	15'h5301: q<=8'h1c;
	15'h5302: q<=8'h38;
	15'h5303: q<=8'h3e;
	15'h5304: q<=8'h1e;
	15'h5305: q<=8'h1a;
	15'h5306: q<=8'h2a;
	15'h5307: q<=8'h1e;
	15'h5308: q<=8'h30;
	15'h5309: q<=8'h00;
	15'h530a: q<=8'h42;
	15'h530b: q<=8'h1e;
	15'h530c: q<=8'h30;
	15'h530d: q<=8'h30;
	15'h530e: q<=8'h00;
	15'h530f: q<=8'h38;
	15'h5310: q<=8'h26;
	15'h5311: q<=8'h1a;
	15'h5312: q<=8'h24;
	15'h5313: q<=8'h3c;
	15'h5314: q<=8'h26;
	15'h5315: q<=8'ha2;
	15'h5316: q<=8'hac;
	15'h5317: q<=8'h32;
	15'h5318: q<=8'h34;
	15'h5319: q<=8'h38;
	15'h531a: q<=8'h26;
	15'h531b: q<=8'h2e;
	15'h531c: q<=8'h16;
	15'h531d: q<=8'h00;
	15'h531e: q<=8'h20;
	15'h531f: q<=8'h26;
	15'h5320: q<=8'h38;
	15'h5321: q<=8'h1e;
	15'h5322: q<=8'h00;
	15'h5323: q<=8'h34;
	15'h5324: q<=8'h16;
	15'h5325: q<=8'h38;
	15'h5326: q<=8'h16;
	15'h5327: q<=8'h00;
	15'h5328: q<=8'h3a;
	15'h5329: q<=8'h1e;
	15'h532a: q<=8'h2c;
	15'h532b: q<=8'h1e;
	15'h532c: q<=8'h1a;
	15'h532d: q<=8'h1a;
	15'h532e: q<=8'h26;
	15'h532f: q<=8'h32;
	15'h5330: q<=8'h30;
	15'h5331: q<=8'h16;
	15'h5332: q<=8'hb8;
	15'h5333: q<=8'hbc;
	15'h5334: q<=8'h24;
	15'h5335: q<=8'h26;
	15'h5336: q<=8'h22;
	15'h5337: q<=8'h24;
	15'h5338: q<=8'h00;
	15'h5339: q<=8'h3a;
	15'h533a: q<=8'h1a;
	15'h533b: q<=8'h32;
	15'h533c: q<=8'h38;
	15'h533d: q<=8'h1e;
	15'h533e: q<=8'hba;
	15'h533f: q<=8'h9e;
	15'h5340: q<=8'h2e;
	15'h5341: q<=8'h1e;
	15'h5342: q<=8'h26;
	15'h5343: q<=8'h2c;
	15'h5344: q<=8'h2c;
	15'h5345: q<=8'h1e;
	15'h5346: q<=8'h3e;
	15'h5347: q<=8'h38;
	15'h5348: q<=8'h3a;
	15'h5349: q<=8'h00;
	15'h534a: q<=8'h3a;
	15'h534b: q<=8'h1a;
	15'h534c: q<=8'h32;
	15'h534d: q<=8'h38;
	15'h534e: q<=8'h1e;
	15'h534f: q<=8'hba;
	15'h5350: q<=8'hb0;
	15'h5351: q<=8'h24;
	15'h5352: q<=8'h32;
	15'h5353: q<=8'h1e;
	15'h5354: q<=8'h1a;
	15'h5355: q<=8'h24;
	15'h5356: q<=8'h3a;
	15'h5357: q<=8'h3c;
	15'h5358: q<=8'h48;
	15'h5359: q<=8'h16;
	15'h535a: q<=8'h24;
	15'h535b: q<=8'h2c;
	15'h535c: q<=8'h1e;
	15'h535d: q<=8'hb0;
	15'h535e: q<=8'hd4;
	15'h535f: q<=8'h38;
	15'h5360: q<=8'h1e;
	15'h5361: q<=8'h1a;
	15'h5362: q<=8'h32;
	15'h5363: q<=8'h38;
	15'h5364: q<=8'h1c;
	15'h5365: q<=8'hba;
	15'h5366: q<=8'hc2;
	15'h5367: q<=8'h38;
	15'h5368: q<=8'h16;
	15'h5369: q<=8'h30;
	15'h536a: q<=8'h2a;
	15'h536b: q<=8'h26;
	15'h536c: q<=8'h30;
	15'h536d: q<=8'h22;
	15'h536e: q<=8'h00;
	15'h536f: q<=8'h20;
	15'h5370: q<=8'h38;
	15'h5371: q<=8'h32;
	15'h5372: q<=8'h2e;
	15'h5373: q<=8'h00;
	15'h5374: q<=8'h04;
	15'h5375: q<=8'h00;
	15'h5376: q<=8'h3c;
	15'h5377: q<=8'h32;
	15'h5378: q<=8'h80;
	15'h5379: q<=8'hc2;
	15'h537a: q<=8'h34;
	15'h537b: q<=8'h2c;
	15'h537c: q<=8'h16;
	15'h537d: q<=8'h1a;
	15'h537e: q<=8'h1e;
	15'h537f: q<=8'h2e;
	15'h5380: q<=8'h1e;
	15'h5381: q<=8'h30;
	15'h5382: q<=8'h3c;
	15'h5383: q<=8'h00;
	15'h5384: q<=8'h1c;
	15'h5385: q<=8'h1e;
	15'h5386: q<=8'h00;
	15'h5387: q<=8'h04;
	15'h5388: q<=8'h00;
	15'h5389: q<=8'h16;
	15'h538a: q<=8'h80;
	15'h538b: q<=8'hbc;
	15'h538c: q<=8'h38;
	15'h538d: q<=8'h16;
	15'h538e: q<=8'h30;
	15'h538f: q<=8'h22;
	15'h5390: q<=8'h2c;
	15'h5391: q<=8'h26;
	15'h5392: q<=8'h3a;
	15'h5393: q<=8'h3c;
	15'h5394: q<=8'h1e;
	15'h5395: q<=8'h00;
	15'h5396: q<=8'h40;
	15'h5397: q<=8'h32;
	15'h5398: q<=8'h30;
	15'h5399: q<=8'h00;
	15'h539a: q<=8'h04;
	15'h539b: q<=8'h00;
	15'h539c: q<=8'h48;
	15'h539d: q<=8'h3e;
	15'h539e: q<=8'h2e;
	15'h539f: q<=8'h80;
	15'h53a0: q<=8'hc8;
	15'h53a1: q<=8'h38;
	15'h53a2: q<=8'h16;
	15'h53a3: q<=8'h30;
	15'h53a4: q<=8'h2a;
	15'h53a5: q<=8'h26;
	15'h53a6: q<=8'h30;
	15'h53a7: q<=8'h22;
	15'h53a8: q<=8'h00;
	15'h53a9: q<=8'h1c;
	15'h53aa: q<=8'h1e;
	15'h53ab: q<=8'h00;
	15'h53ac: q<=8'h04;
	15'h53ad: q<=8'h00;
	15'h53ae: q<=8'h16;
	15'h53af: q<=8'h80;
	15'h53b0: q<=8'hd9;
	15'h53b1: q<=8'h38;
	15'h53b2: q<=8'h16;
	15'h53b3: q<=8'h3c;
	15'h53b4: q<=8'h1e;
	15'h53b5: q<=8'h00;
	15'h53b6: q<=8'h46;
	15'h53b7: q<=8'h32;
	15'h53b8: q<=8'h3e;
	15'h53b9: q<=8'h38;
	15'h53ba: q<=8'h3a;
	15'h53bb: q<=8'h1e;
	15'h53bc: q<=8'h2c;
	15'h53bd: q<=8'ha0;
	15'h53be: q<=8'hdc;
	15'h53bf: q<=8'h1e;
	15'h53c0: q<=8'h40;
	15'h53c1: q<=8'h16;
	15'h53c2: q<=8'h2c;
	15'h53c3: q<=8'h3e;
	15'h53c4: q<=8'h1e;
	15'h53c5: q<=8'h48;
	15'h53c6: q<=8'h4c;
	15'h53c7: q<=8'h40;
	15'h53c8: q<=8'h32;
	15'h53c9: q<=8'h3e;
	15'h53ca: q<=8'hba;
	15'h53cb: q<=8'hd6;
	15'h53cc: q<=8'h3a;
	15'h53cd: q<=8'h1e;
	15'h53ce: q<=8'h2c;
	15'h53cf: q<=8'h18;
	15'h53d0: q<=8'h3a;
	15'h53d1: q<=8'h3c;
	15'h53d2: q<=8'h00;
	15'h53d3: q<=8'h38;
	15'h53d4: q<=8'h1e;
	15'h53d5: q<=8'h1a;
	15'h53d6: q<=8'h24;
	15'h53d7: q<=8'h30;
	15'h53d8: q<=8'h1e;
	15'h53d9: q<=8'hb0;
	15'h53da: q<=8'hdf;
	15'h53db: q<=8'h1a;
	15'h53dc: q<=8'h16;
	15'h53dd: q<=8'h2c;
	15'h53de: q<=8'h26;
	15'h53df: q<=8'h20;
	15'h53e0: q<=8'h26;
	15'h53e1: q<=8'h36;
	15'h53e2: q<=8'h3e;
	15'h53e3: q<=8'h1e;
	15'h53e4: q<=8'h3a;
	15'h53e5: q<=8'h9e;
	15'h53e6: q<=8'haa;
	15'h53e7: q<=8'h30;
	15'h53e8: q<=8'h32;
	15'h53e9: q<=8'h40;
	15'h53ea: q<=8'h26;
	15'h53eb: q<=8'h1a;
	15'h53ec: q<=8'h9e;
	15'h53ed: q<=8'haa;
	15'h53ee: q<=8'h30;
	15'h53ef: q<=8'h32;
	15'h53f0: q<=8'h40;
	15'h53f1: q<=8'h26;
	15'h53f2: q<=8'h1a;
	15'h53f3: q<=8'h26;
	15'h53f4: q<=8'hb2;
	15'h53f5: q<=8'haa;
	15'h53f6: q<=8'h16;
	15'h53f7: q<=8'h30;
	15'h53f8: q<=8'h20;
	15'h53f9: q<=8'h16;
	15'h53fa: q<=8'h1e;
	15'h53fb: q<=8'h30;
	15'h53fc: q<=8'h22;
	15'h53fd: q<=8'h1e;
	15'h53fe: q<=8'hb8;
	15'h53ff: q<=8'h4a;
	15'h5400: q<=8'h1e;
	15'h5401: q<=8'h44;
	15'h5402: q<=8'h34;
	15'h5403: q<=8'h1e;
	15'h5404: q<=8'h38;
	15'h5405: q<=8'hbc;
	15'h5406: q<=8'h45;
	15'h5407: q<=8'h1e;
	15'h5408: q<=8'h44;
	15'h5409: q<=8'h34;
	15'h540a: q<=8'h1e;
	15'h540b: q<=8'h38;
	15'h540c: q<=8'h3c;
	15'h540d: q<=8'hb2;
	15'h540e: q<=8'h40;
	15'h540f: q<=8'h1e;
	15'h5410: q<=8'h38;
	15'h5411: q<=8'h20;
	15'h5412: q<=8'h16;
	15'h5413: q<=8'h24;
	15'h5414: q<=8'h38;
	15'h5415: q<=8'h1e;
	15'h5416: q<=8'hb0;
	15'h5417: q<=8'h8b;
	15'h5418: q<=8'h18;
	15'h5419: q<=8'h32;
	15'h541a: q<=8'h30;
	15'h541b: q<=8'h3e;
	15'h541c: q<=8'hba;
	15'h541d: q<=8'he8;
	15'h541e: q<=8'h3c;
	15'h541f: q<=8'h26;
	15'h5420: q<=8'h2e;
	15'h5421: q<=8'h9e;
	15'h5422: q<=8'he0;
	15'h5423: q<=8'h1c;
	15'h5424: q<=8'h3e;
	15'h5425: q<=8'h38;
	15'h5426: q<=8'h1e;
	15'h5427: q<=8'h9e;
	15'h5428: q<=8'he8;
	15'h5429: q<=8'h48;
	15'h542a: q<=8'h1e;
	15'h542b: q<=8'h26;
	15'h542c: q<=8'hbc;
	15'h542d: q<=8'he4;
	15'h542e: q<=8'h3c;
	15'h542f: q<=8'h26;
	15'h5430: q<=8'h1e;
	15'h5431: q<=8'h2e;
	15'h5432: q<=8'h34;
	15'h5433: q<=8'hb2;
	15'h5434: q<=8'h8b;
	15'h5435: q<=8'h2c;
	15'h5436: q<=8'h1e;
	15'h5437: q<=8'h40;
	15'h5438: q<=8'h1e;
	15'h5439: q<=8'hac;
	15'h543a: q<=8'h8b;
	15'h543b: q<=8'h30;
	15'h543c: q<=8'h26;
	15'h543d: q<=8'h40;
	15'h543e: q<=8'h1e;
	15'h543f: q<=8'h16;
	15'h5440: q<=8'hbe;
	15'h5441: q<=8'h8b;
	15'h5442: q<=8'h22;
	15'h5443: q<=8'h38;
	15'h5444: q<=8'h16;
	15'h5445: q<=8'h9c;
	15'h5446: q<=8'h8b;
	15'h5447: q<=8'h30;
	15'h5448: q<=8'h26;
	15'h5449: q<=8'h40;
	15'h544a: q<=8'h1e;
	15'h544b: q<=8'hac;
	15'h544c: q<=8'h8b;
	15'h544d: q<=8'h24;
	15'h544e: q<=8'h32;
	15'h544f: q<=8'h2c;
	15'h5450: q<=8'h9e;
	15'h5451: q<=8'h8b;
	15'h5452: q<=8'h3c;
	15'h5453: q<=8'h38;
	15'h5454: q<=8'h32;
	15'h5455: q<=8'hbe;
	15'h5456: q<=8'h8b;
	15'h5457: q<=8'h24;
	15'h5458: q<=8'h32;
	15'h5459: q<=8'h46;
	15'h545a: q<=8'hb2;
	15'h545b: q<=8'h8b;
	15'h545c: q<=8'h2c;
	15'h545d: q<=8'h32;
	15'h545e: q<=8'h1a;
	15'h545f: q<=8'ha4;
	15'h5460: q<=8'hdc;
	15'h5461: q<=8'h26;
	15'h5462: q<=8'h30;
	15'h5463: q<=8'h3a;
	15'h5464: q<=8'h1e;
	15'h5465: q<=8'h38;
	15'h5466: q<=8'h3c;
	15'h5467: q<=8'h00;
	15'h5468: q<=8'h1a;
	15'h5469: q<=8'h32;
	15'h546a: q<=8'h26;
	15'h546b: q<=8'h30;
	15'h546c: q<=8'hba;
	15'h546d: q<=8'hc1;
	15'h546e: q<=8'h26;
	15'h546f: q<=8'h30;
	15'h5470: q<=8'h3c;
	15'h5471: q<=8'h38;
	15'h5472: q<=8'h32;
	15'h5473: q<=8'h1c;
	15'h5474: q<=8'h3e;
	15'h5475: q<=8'h26;
	15'h5476: q<=8'h38;
	15'h5477: q<=8'h1e;
	15'h5478: q<=8'h00;
	15'h5479: q<=8'h2c;
	15'h547a: q<=8'h1e;
	15'h547b: q<=8'h3a;
	15'h547c: q<=8'h00;
	15'h547d: q<=8'h34;
	15'h547e: q<=8'h26;
	15'h547f: q<=8'h1e;
	15'h5480: q<=8'h1a;
	15'h5481: q<=8'h1e;
	15'h5482: q<=8'hba;
	15'h5483: q<=8'hd6;
	15'h5484: q<=8'h22;
	15'h5485: q<=8'h1e;
	15'h5486: q<=8'h2c;
	15'h5487: q<=8'h1c;
	15'h5488: q<=8'h00;
	15'h5489: q<=8'h1e;
	15'h548a: q<=8'h26;
	15'h548b: q<=8'h30;
	15'h548c: q<=8'h42;
	15'h548d: q<=8'h1e;
	15'h548e: q<=8'h38;
	15'h548f: q<=8'h20;
	15'h5490: q<=8'h1e;
	15'h5491: q<=8'hb0;
	15'h5492: q<=8'hd6;
	15'h5493: q<=8'h26;
	15'h5494: q<=8'h30;
	15'h5495: q<=8'h3a;
	15'h5496: q<=8'h1e;
	15'h5497: q<=8'h38;
	15'h5498: q<=8'h3c;
	15'h5499: q<=8'h1e;
	15'h549a: q<=8'h00;
	15'h549b: q<=8'h20;
	15'h549c: q<=8'h26;
	15'h549d: q<=8'h1a;
	15'h549e: q<=8'h24;
	15'h549f: q<=8'h16;
	15'h54a0: q<=8'hba;
	15'h54a1: q<=8'h00;
	15'h54a2: q<=8'h20;
	15'h54a3: q<=8'h38;
	15'h54a4: q<=8'h1e;
	15'h54a5: q<=8'h1e;
	15'h54a6: q<=8'h00;
	15'h54a7: q<=8'h34;
	15'h54a8: q<=8'h2c;
	15'h54a9: q<=8'h16;
	15'h54aa: q<=8'hc6;
	15'h54ab: q<=8'h0e;
	15'h54ac: q<=8'h04;
	15'h54ad: q<=8'h00;
	15'h54ae: q<=8'h1a;
	15'h54af: q<=8'h32;
	15'h54b0: q<=8'h26;
	15'h54b1: q<=8'h30;
	15'h54b2: q<=8'h00;
	15'h54b3: q<=8'h06;
	15'h54b4: q<=8'h00;
	15'h54b5: q<=8'h34;
	15'h54b6: q<=8'h2c;
	15'h54b7: q<=8'h16;
	15'h54b8: q<=8'h46;
	15'h54b9: q<=8'hba;
	15'h54ba: q<=8'hfa;
	15'h54bb: q<=8'h04;
	15'h54bc: q<=8'h00;
	15'h54bd: q<=8'h34;
	15'h54be: q<=8'h26;
	15'h54bf: q<=8'h1e;
	15'h54c0: q<=8'h1a;
	15'h54c1: q<=8'h1e;
	15'h54c2: q<=8'h00;
	15'h54c3: q<=8'h06;
	15'h54c4: q<=8'h00;
	15'h54c5: q<=8'h28;
	15'h54c6: q<=8'h32;
	15'h54c7: q<=8'h3e;
	15'h54c8: q<=8'h1e;
	15'h54c9: q<=8'h3e;
	15'h54ca: q<=8'h38;
	15'h54cb: q<=8'hba;
	15'h54cc: q<=8'h00;
	15'h54cd: q<=8'h04;
	15'h54ce: q<=8'h00;
	15'h54cf: q<=8'h2e;
	15'h54d0: q<=8'h3e;
	15'h54d1: q<=8'h1e;
	15'h54d2: q<=8'h30;
	15'h54d3: q<=8'h48;
	15'h54d4: q<=8'h00;
	15'h54d5: q<=8'h06;
	15'h54d6: q<=8'h00;
	15'h54d7: q<=8'h3a;
	15'h54d8: q<=8'h34;
	15'h54d9: q<=8'h26;
	15'h54da: q<=8'h1e;
	15'h54db: q<=8'h2c;
	15'h54dc: q<=8'h9e;
	15'h54dd: q<=8'hfa;
	15'h54de: q<=8'h04;
	15'h54df: q<=8'h00;
	15'h54e0: q<=8'h2e;
	15'h54e1: q<=8'h32;
	15'h54e2: q<=8'h30;
	15'h54e3: q<=8'h1e;
	15'h54e4: q<=8'h1c;
	15'h54e5: q<=8'h16;
	15'h54e6: q<=8'h00;
	15'h54e7: q<=8'h06;
	15'h54e8: q<=8'h00;
	15'h54e9: q<=8'h28;
	15'h54ea: q<=8'h3e;
	15'h54eb: q<=8'h1e;
	15'h54ec: q<=8'h22;
	15'h54ed: q<=8'h32;
	15'h54ee: q<=8'hba;
	15'h54ef: q<=8'h14;
	15'h54f0: q<=8'h04;
	15'h54f1: q<=8'h00;
	15'h54f2: q<=8'h1a;
	15'h54f3: q<=8'h32;
	15'h54f4: q<=8'h26;
	15'h54f5: q<=8'h30;
	15'h54f6: q<=8'h00;
	15'h54f7: q<=8'h04;
	15'h54f8: q<=8'h00;
	15'h54f9: q<=8'h34;
	15'h54fa: q<=8'h2c;
	15'h54fb: q<=8'h16;
	15'h54fc: q<=8'hc6;
	15'h54fd: q<=8'h00;
	15'h54fe: q<=8'h04;
	15'h54ff: q<=8'h00;
	15'h5500: q<=8'h34;
	15'h5501: q<=8'h26;
	15'h5502: q<=8'h1e;
	15'h5503: q<=8'h1a;
	15'h5504: q<=8'h1e;
	15'h5505: q<=8'h00;
	15'h5506: q<=8'h04;
	15'h5507: q<=8'h00;
	15'h5508: q<=8'h28;
	15'h5509: q<=8'h32;
	15'h550a: q<=8'h3e;
	15'h550b: q<=8'h1e;
	15'h550c: q<=8'h3e;
	15'h550d: q<=8'hb8;
	15'h550e: q<=8'h00;
	15'h550f: q<=8'h04;
	15'h5510: q<=8'h00;
	15'h5511: q<=8'h2e;
	15'h5512: q<=8'h3e;
	15'h5513: q<=8'h1e;
	15'h5514: q<=8'h30;
	15'h5515: q<=8'h48;
	15'h5516: q<=8'h1e;
	15'h5517: q<=8'h00;
	15'h5518: q<=8'h04;
	15'h5519: q<=8'h00;
	15'h551a: q<=8'h3a;
	15'h551b: q<=8'h34;
	15'h551c: q<=8'h26;
	15'h551d: q<=8'h1e;
	15'h551e: q<=8'hac;
	15'h551f: q<=8'h00;
	15'h5520: q<=8'h04;
	15'h5521: q<=8'h00;
	15'h5522: q<=8'h2e;
	15'h5523: q<=8'h32;
	15'h5524: q<=8'h30;
	15'h5525: q<=8'h1e;
	15'h5526: q<=8'h1c;
	15'h5527: q<=8'h16;
	15'h5528: q<=8'h00;
	15'h5529: q<=8'h04;
	15'h552a: q<=8'h00;
	15'h552b: q<=8'h28;
	15'h552c: q<=8'h3e;
	15'h552d: q<=8'h1e;
	15'h552e: q<=8'h22;
	15'h552f: q<=8'hb2;
	15'h5530: q<=8'h0e;
	15'h5531: q<=8'h06;
	15'h5532: q<=8'h00;
	15'h5533: q<=8'h1a;
	15'h5534: q<=8'h32;
	15'h5535: q<=8'h26;
	15'h5536: q<=8'h30;
	15'h5537: q<=8'h3a;
	15'h5538: q<=8'h00;
	15'h5539: q<=8'h04;
	15'h553a: q<=8'h00;
	15'h553b: q<=8'h34;
	15'h553c: q<=8'h2c;
	15'h553d: q<=8'h16;
	15'h553e: q<=8'hc6;
	15'h553f: q<=8'hfa;
	15'h5540: q<=8'h06;
	15'h5541: q<=8'h00;
	15'h5542: q<=8'h34;
	15'h5543: q<=8'h26;
	15'h5544: q<=8'h1e;
	15'h5545: q<=8'h1a;
	15'h5546: q<=8'h1e;
	15'h5547: q<=8'h3a;
	15'h5548: q<=8'h00;
	15'h5549: q<=8'h04;
	15'h554a: q<=8'h00;
	15'h554b: q<=8'h28;
	15'h554c: q<=8'h32;
	15'h554d: q<=8'h3e;
	15'h554e: q<=8'h1e;
	15'h554f: q<=8'h3e;
	15'h5550: q<=8'hb8;
	15'h5551: q<=8'hfa;
	15'h5552: q<=8'h06;
	15'h5553: q<=8'h00;
	15'h5554: q<=8'h2e;
	15'h5555: q<=8'h3e;
	15'h5556: q<=8'h1e;
	15'h5557: q<=8'h30;
	15'h5558: q<=8'h48;
	15'h5559: q<=8'h1e;
	15'h555a: q<=8'h30;
	15'h555b: q<=8'h00;
	15'h555c: q<=8'h04;
	15'h555d: q<=8'h00;
	15'h555e: q<=8'h3a;
	15'h555f: q<=8'h34;
	15'h5560: q<=8'h26;
	15'h5561: q<=8'h1e;
	15'h5562: q<=8'hac;
	15'h5563: q<=8'hfa;
	15'h5564: q<=8'h06;
	15'h5565: q<=8'h00;
	15'h5566: q<=8'h2e;
	15'h5567: q<=8'h32;
	15'h5568: q<=8'h30;
	15'h5569: q<=8'h1e;
	15'h556a: q<=8'h1c;
	15'h556b: q<=8'h16;
	15'h556c: q<=8'h3a;
	15'h556d: q<=8'h00;
	15'h556e: q<=8'h04;
	15'h556f: q<=8'h00;
	15'h5570: q<=8'h28;
	15'h5571: q<=8'h3e;
	15'h5572: q<=8'h1e;
	15'h5573: q<=8'h22;
	15'h5574: q<=8'hb2;
	15'h5575: q<=8'hd3;
	15'h5576: q<=8'h50;
	15'h5577: q<=8'h00;
	15'h5578: q<=8'h2e;
	15'h5579: q<=8'h1a;
	15'h557a: q<=8'h2e;
	15'h557b: q<=8'h2c;
	15'h557c: q<=8'h44;
	15'h557d: q<=8'h44;
	15'h557e: q<=8'h44;
	15'h557f: q<=8'h00;
	15'h5580: q<=8'h16;
	15'h5581: q<=8'h3c;
	15'h5582: q<=8'h16;
	15'h5583: q<=8'h38;
	15'h5584: q<=8'ha6;
	15'h5585: q<=8'ha0;
	15'h5586: q<=8'h1a;
	15'h5587: q<=8'h38;
	15'h5588: q<=8'h1e;
	15'h5589: q<=8'h1c;
	15'h558a: q<=8'h26;
	15'h558b: q<=8'h3c;
	15'h558c: q<=8'h3a;
	15'h558d: q<=8'h80;
	15'h558e: q<=8'ha0;
	15'h558f: q<=8'h2a;
	15'h5590: q<=8'h38;
	15'h5591: q<=8'h1e;
	15'h5592: q<=8'h1c;
	15'h5593: q<=8'h26;
	15'h5594: q<=8'h3c;
	15'h5595: q<=8'h1e;
	15'h5596: q<=8'h80;
	15'h5597: q<=8'ha0;
	15'h5598: q<=8'h1a;
	15'h5599: q<=8'h38;
	15'h559a: q<=8'h1e;
	15'h559b: q<=8'h1c;
	15'h559c: q<=8'h26;
	15'h559d: q<=8'h3c;
	15'h559e: q<=8'h32;
	15'h559f: q<=8'h3a;
	15'h55a0: q<=8'h80;
	15'h55a1: q<=8'hda;
	15'h55a2: q<=8'h18;
	15'h55a3: q<=8'h32;
	15'h55a4: q<=8'h30;
	15'h55a5: q<=8'h3e;
	15'h55a6: q<=8'h3a;
	15'h55a7: q<=8'h80;
	15'h55a8: q<=8'hd0;
	15'h55a9: q<=8'h06;
	15'h55aa: q<=8'h00;
	15'h55ab: q<=8'h1a;
	15'h55ac: q<=8'h38;
	15'h55ad: q<=8'h1e;
	15'h55ae: q<=8'h1c;
	15'h55af: q<=8'h26;
	15'h55b0: q<=8'h3c;
	15'h55b1: q<=8'h00;
	15'h55b2: q<=8'h2e;
	15'h55b3: q<=8'h26;
	15'h55b4: q<=8'h30;
	15'h55b5: q<=8'h26;
	15'h55b6: q<=8'h2e;
	15'h55b7: q<=8'h3e;
	15'h55b8: q<=8'hae;
	15'h55b9: q<=8'hd6;
	15'h55ba: q<=8'h06;
	15'h55bb: q<=8'h00;
	15'h55bc: q<=8'h28;
	15'h55bd: q<=8'h1e;
	15'h55be: q<=8'h3e;
	15'h55bf: q<=8'h44;
	15'h55c0: q<=8'h00;
	15'h55c1: q<=8'h2e;
	15'h55c2: q<=8'h26;
	15'h55c3: q<=8'h30;
	15'h55c4: q<=8'h26;
	15'h55c5: q<=8'h2e;
	15'h55c6: q<=8'h3e;
	15'h55c7: q<=8'hae;
	15'h55c8: q<=8'hd0;
	15'h55c9: q<=8'h06;
	15'h55ca: q<=8'h00;
	15'h55cb: q<=8'h3a;
	15'h55cc: q<=8'h34;
	15'h55cd: q<=8'h26;
	15'h55ce: q<=8'h1e;
	15'h55cf: q<=8'h2c;
	15'h55d0: q<=8'h1e;
	15'h55d1: q<=8'h00;
	15'h55d2: q<=8'h2e;
	15'h55d3: q<=8'h26;
	15'h55d4: q<=8'h30;
	15'h55d5: q<=8'h26;
	15'h55d6: q<=8'h2e;
	15'h55d7: q<=8'h3e;
	15'h55d8: q<=8'hae;
	15'h55d9: q<=8'hd3;
	15'h55da: q<=8'h06;
	15'h55db: q<=8'h00;
	15'h55dc: q<=8'h28;
	15'h55dd: q<=8'h3e;
	15'h55de: q<=8'h1e;
	15'h55df: q<=8'h22;
	15'h55e0: q<=8'h32;
	15'h55e1: q<=8'h3a;
	15'h55e2: q<=8'h00;
	15'h55e3: q<=8'h2e;
	15'h55e4: q<=8'h26;
	15'h55e5: q<=8'h30;
	15'h55e6: q<=8'h26;
	15'h55e7: q<=8'h2e;
	15'h55e8: q<=8'hb2;
	15'h55e9: q<=8'hc8;
	15'h55ea: q<=8'h18;
	15'h55eb: q<=8'h32;
	15'h55ec: q<=8'h30;
	15'h55ed: q<=8'h3e;
	15'h55ee: q<=8'h3a;
	15'h55ef: q<=8'h00;
	15'h55f0: q<=8'h1e;
	15'h55f1: q<=8'h40;
	15'h55f2: q<=8'h1e;
	15'h55f3: q<=8'h38;
	15'h55f4: q<=8'h46;
	15'h55f5: q<=8'h80;
	15'h55f6: q<=8'hce;
	15'h55f7: q<=8'h18;
	15'h55f8: q<=8'h32;
	15'h55f9: q<=8'h30;
	15'h55fa: q<=8'h3e;
	15'h55fb: q<=8'h3a;
	15'h55fc: q<=8'h00;
	15'h55fd: q<=8'h1a;
	15'h55fe: q<=8'h24;
	15'h55ff: q<=8'h16;
	15'h5600: q<=8'h36;
	15'h5601: q<=8'h3e;
	15'h5602: q<=8'h1e;
	15'h5603: q<=8'h80;
	15'h5604: q<=8'hce;
	15'h5605: q<=8'h18;
	15'h5606: q<=8'h32;
	15'h5607: q<=8'h30;
	15'h5608: q<=8'h3e;
	15'h5609: q<=8'h3a;
	15'h560a: q<=8'h00;
	15'h560b: q<=8'h28;
	15'h560c: q<=8'h1e;
	15'h560d: q<=8'h1c;
	15'h560e: q<=8'h1e;
	15'h560f: q<=8'h80;
	15'h5610: q<=8'hc8;
	15'h5611: q<=8'h18;
	15'h5612: q<=8'h32;
	15'h5613: q<=8'h30;
	15'h5614: q<=8'h3e;
	15'h5615: q<=8'h3a;
	15'h5616: q<=8'h00;
	15'h5617: q<=8'h1a;
	15'h5618: q<=8'h16;
	15'h5619: q<=8'h1c;
	15'h561a: q<=8'h16;
	15'h561b: q<=8'h80;
	15'h561c: q<=8'hb8;
	15'h561d: q<=8'h16;
	15'h561e: q<=8'h40;
	15'h561f: q<=8'h32;
	15'h5620: q<=8'h26;
	15'h5621: q<=8'h1c;
	15'h5622: q<=8'h00;
	15'h5623: q<=8'h3a;
	15'h5624: q<=8'h34;
	15'h5625: q<=8'h26;
	15'h5626: q<=8'h2a;
	15'h5627: q<=8'h1e;
	15'h5628: q<=8'hba;
	15'h5629: q<=8'h88;
	15'h562a: q<=8'h16;
	15'h562b: q<=8'h3c;
	15'h562c: q<=8'h3c;
	15'h562d: q<=8'h1e;
	15'h562e: q<=8'h30;
	15'h562f: q<=8'h3c;
	15'h5630: q<=8'h26;
	15'h5631: q<=8'h32;
	15'h5632: q<=8'h30;
	15'h5633: q<=8'h00;
	15'h5634: q<=8'h16;
	15'h5635: q<=8'h3e;
	15'h5636: q<=8'h44;
	15'h5637: q<=8'h00;
	15'h5638: q<=8'h2c;
	15'h5639: q<=8'h16;
	15'h563a: q<=8'h30;
	15'h563b: q<=8'h1a;
	15'h563c: q<=8'h1e;
	15'h563d: q<=8'hba;
	15'h563e: q<=8'h96;
	15'h563f: q<=8'h3a;
	15'h5640: q<=8'h34;
	15'h5641: q<=8'h26;
	15'h5642: q<=8'h3c;
	15'h5643: q<=8'h48;
	15'h5644: q<=8'h1e;
	15'h5645: q<=8'h30;
	15'h5646: q<=8'h00;
	15'h5647: q<=8'h16;
	15'h5648: q<=8'h3e;
	15'h5649: q<=8'h3a;
	15'h564a: q<=8'h42;
	15'h564b: q<=8'h1e;
	15'h564c: q<=8'h26;
	15'h564d: q<=8'h1a;
	15'h564e: q<=8'h24;
	15'h564f: q<=8'h1e;
	15'h5650: q<=8'hb0;
	15'h5651: q<=8'ha0;
	15'h5652: q<=8'h1e;
	15'h5653: q<=8'h40;
	15'h5654: q<=8'h26;
	15'h5655: q<=8'h3c;
	15'h5656: q<=8'h1e;
	15'h5657: q<=8'h00;
	15'h5658: q<=8'h2c;
	15'h5659: q<=8'h16;
	15'h565a: q<=8'h3a;
	15'h565b: q<=8'h00;
	15'h565c: q<=8'h34;
	15'h565d: q<=8'h3e;
	15'h565e: q<=8'h30;
	15'h565f: q<=8'h3c;
	15'h5660: q<=8'h16;
	15'h5661: q<=8'hba;
	15'h5662: q<=8'he0;
	15'h5663: q<=8'h2c;
	15'h5664: q<=8'h1e;
	15'h5665: q<=8'h40;
	15'h5666: q<=8'h1e;
	15'h5667: q<=8'hac;
	15'h5668: q<=8'hda;
	15'h5669: q<=8'h30;
	15'h566a: q<=8'h26;
	15'h566b: q<=8'h40;
	15'h566c: q<=8'h1e;
	15'h566d: q<=8'h16;
	15'h566e: q<=8'hbe;
	15'h566f: q<=8'he2;
	15'h5670: q<=8'h22;
	15'h5671: q<=8'h38;
	15'h5672: q<=8'h16;
	15'h5673: q<=8'h9c;
	15'h5674: q<=8'he0;
	15'h5675: q<=8'h30;
	15'h5676: q<=8'h26;
	15'h5677: q<=8'h40;
	15'h5678: q<=8'h1e;
	15'h5679: q<=8'hac;
	15'h567a: q<=8'hc4;
	15'h567b: q<=8'h3a;
	15'h567c: q<=8'h3e;
	15'h567d: q<=8'h34;
	15'h567e: q<=8'h1e;
	15'h567f: q<=8'h38;
	15'h5680: q<=8'h48;
	15'h5681: q<=8'h16;
	15'h5682: q<=8'h34;
	15'h5683: q<=8'h34;
	15'h5684: q<=8'h1e;
	15'h5685: q<=8'h38;
	15'h5686: q<=8'h00;
	15'h5687: q<=8'h38;
	15'h5688: q<=8'h1e;
	15'h5689: q<=8'h1a;
	15'h568a: q<=8'h24;
	15'h568b: q<=8'h16;
	15'h568c: q<=8'h38;
	15'h568d: q<=8'h22;
	15'h568e: q<=8'h9e;
	15'h568f: q<=8'hcd;
	15'h5690: q<=8'h30;
	15'h5691: q<=8'h1e;
	15'h5692: q<=8'h3e;
	15'h5693: q<=8'h1e;
	15'h5694: q<=8'h38;
	15'h5695: q<=8'h00;
	15'h5696: q<=8'h3a;
	15'h5697: q<=8'h3e;
	15'h5698: q<=8'h34;
	15'h5699: q<=8'h1e;
	15'h569a: q<=8'h38;
	15'h569b: q<=8'h48;
	15'h569c: q<=8'h16;
	15'h569d: q<=8'h34;
	15'h569e: q<=8'h34;
	15'h569f: q<=8'h1e;
	15'h56a0: q<=8'hb8;
	15'h56a1: q<=8'hcd;
	15'h56a2: q<=8'h30;
	15'h56a3: q<=8'h3e;
	15'h56a4: q<=8'h1e;
	15'h56a5: q<=8'h40;
	15'h56a6: q<=8'h32;
	15'h56a7: q<=8'h00;
	15'h56a8: q<=8'h3a;
	15'h56a9: q<=8'h3e;
	15'h56aa: q<=8'h34;
	15'h56ab: q<=8'h1e;
	15'h56ac: q<=8'h38;
	15'h56ad: q<=8'h48;
	15'h56ae: q<=8'h16;
	15'h56af: q<=8'h34;
	15'h56b0: q<=8'h34;
	15'h56b1: q<=8'h1e;
	15'h56b2: q<=8'hb8;
	15'h56b3: q<=8'h31;
	15'h56b4: q<=8'hd0;
	15'h56b5: q<=8'h6d;
	15'h56b6: q<=8'hd0;
	15'h56b7: q<=8'ha9;
	15'h56b8: q<=8'hd0;
	15'h56b9: q<=8'he5;
	15'h56ba: q<=8'hd0;
	15'h56bb: q<=8'had;
	15'h56bc: q<=8'h00;
	15'h56bd: q<=8'h0e;
	15'h56be: q<=8'h85;
	15'h56bf: q<=8'h0a;
	15'h56c0: q<=8'h29;
	15'h56c1: q<=8'h38;
	15'h56c2: q<=8'h4a;
	15'h56c3: q<=8'h4a;
	15'h56c4: q<=8'h4a;
	15'h56c5: q<=8'haa;
	15'h56c6: q<=8'hbd;
	15'h56c7: q<=8'hf7;
	15'h56c8: q<=8'hd6;
	15'h56c9: q<=8'h8d;
	15'h56ca: q<=8'h56;
	15'h56cb: q<=8'h01;
	15'h56cc: q<=8'had;
	15'h56cd: q<=8'h00;
	15'h56ce: q<=8'h0d;
	15'h56cf: q<=8'h49;
	15'h56d0: q<=8'h02;
	15'h56d1: q<=8'h85;
	15'h56d2: q<=8'h09;
	15'h56d3: q<=8'ha5;
	15'h56d4: q<=8'h0a;
	15'h56d5: q<=8'h2a;
	15'h56d6: q<=8'h2a;
	15'h56d7: q<=8'h2a;
	15'h56d8: q<=8'h29;
	15'h56d9: q<=8'h03;
	15'h56da: q<=8'haa;
	15'h56db: q<=8'hbd;
	15'h56dc: q<=8'hff;
	15'h56dd: q<=8'hd6;
	15'h56de: q<=8'h8d;
	15'h56df: q<=8'h58;
	15'h56e0: q<=8'h01;
	15'h56e1: q<=8'ha5;
	15'h56e2: q<=8'h0a;
	15'h56e3: q<=8'h29;
	15'h56e4: q<=8'h06;
	15'h56e5: q<=8'ha8;
	15'h56e6: q<=8'hb9;
	15'h56e7: q<=8'hb3;
	15'h56e8: q<=8'hd6;
	15'h56e9: q<=8'h85;
	15'h56ea: q<=8'hac;
	15'h56eb: q<=8'hb9;
	15'h56ec: q<=8'hb4;
	15'h56ed: q<=8'hd6;
	15'h56ee: q<=8'h85;
	15'h56ef: q<=8'had;
	15'h56f0: q<=8'h20;
	15'h56f1: q<=8'he0;
	15'h56f2: q<=8'hdb;
	15'h56f3: q<=8'h8d;
	15'h56f4: q<=8'h6a;
	15'h56f5: q<=8'h01;
	15'h56f6: q<=8'h60;
	15'h56f7: q<=8'h02;
	15'h56f8: q<=8'h01;
	15'h56f9: q<=8'h03;
	15'h56fa: q<=8'h04;
	15'h56fb: q<=8'h05;
	15'h56fc: q<=8'h06;
	15'h56fd: q<=8'h07;
	15'h56fe: q<=8'h00;
	15'h56ff: q<=8'h03;
	15'h5700: q<=8'h04;
	15'h5701: q<=8'h05;
	15'h5702: q<=8'h02;
	15'h5703: q<=8'h7c;
	15'h5704: q<=8'h48;
	15'h5705: q<=8'h8a;
	15'h5706: q<=8'h48;
	15'h5707: q<=8'h98;
	15'h5708: q<=8'h48;
	15'h5709: q<=8'hd8;
	15'h570a: q<=8'hba;
	15'h570b: q<=8'he0;
	15'h570c: q<=8'hd0;
	15'h570d: q<=8'h90;
	15'h570e: q<=8'h04;
	15'h570f: q<=8'ha5;
	15'h5710: q<=8'h53;
	15'h5711: q<=8'h10;
	15'h5712: q<=8'h04;
	15'h5713: q<=8'h00;
	15'h5714: q<=8'h4c;
	15'h5715: q<=8'h3f;
	15'h5716: q<=8'hd9;
	15'h5717: q<=8'h8d;
	15'h5718: q<=8'h00;
	15'h5719: q<=8'h50;
	15'h571a: q<=8'h8d;
	15'h571b: q<=8'hcb;
	15'h571c: q<=8'h60;
	15'h571d: q<=8'had;
	15'h571e: q<=8'hc8;
	15'h571f: q<=8'h60;
	15'h5720: q<=8'h49;
	15'h5721: q<=8'h0f;
	15'h5722: q<=8'ha8;
	15'h5723: q<=8'h29;
	15'h5724: q<=8'h10;
	15'h5725: q<=8'h8d;
	15'h5726: q<=8'h17;
	15'h5727: q<=8'h01;
	15'h5728: q<=8'h98;
	15'h5729: q<=8'h38;
	15'h572a: q<=8'he5;
	15'h572b: q<=8'h52;
	15'h572c: q<=8'h29;
	15'h572d: q<=8'h0f;
	15'h572e: q<=8'hc9;
	15'h572f: q<=8'h08;
	15'h5730: q<=8'h90;
	15'h5731: q<=8'h02;
	15'h5732: q<=8'h09;
	15'h5733: q<=8'hf0;
	15'h5734: q<=8'h18;
	15'h5735: q<=8'h65;
	15'h5736: q<=8'h50;
	15'h5737: q<=8'h85;
	15'h5738: q<=8'h50;
	15'h5739: q<=8'h84;
	15'h573a: q<=8'h52;
	15'h573b: q<=8'h8d;
	15'h573c: q<=8'hdb;
	15'h573d: q<=8'h60;
	15'h573e: q<=8'hac;
	15'h573f: q<=8'hd8;
	15'h5740: q<=8'h60;
	15'h5741: q<=8'had;
	15'h5742: q<=8'h00;
	15'h5743: q<=8'h0c;
	15'h5744: q<=8'h85;
	15'h5745: q<=8'h08;
	15'h5746: q<=8'ha5;
	15'h5747: q<=8'h4c;
	15'h5748: q<=8'h84;
	15'h5749: q<=8'h4c;
	15'h574a: q<=8'ha8;
	15'h574b: q<=8'h25;
	15'h574c: q<=8'h4c;
	15'h574d: q<=8'h05;
	15'h574e: q<=8'h4d;
	15'h574f: q<=8'h85;
	15'h5750: q<=8'h4d;
	15'h5751: q<=8'h98;
	15'h5752: q<=8'h05;
	15'h5753: q<=8'h4c;
	15'h5754: q<=8'h25;
	15'h5755: q<=8'h4d;
	15'h5756: q<=8'h85;
	15'h5757: q<=8'h4d;
	15'h5758: q<=8'ha8;
	15'h5759: q<=8'h45;
	15'h575a: q<=8'h4f;
	15'h575b: q<=8'h25;
	15'h575c: q<=8'h4d;
	15'h575d: q<=8'h05;
	15'h575e: q<=8'h4e;
	15'h575f: q<=8'h85;
	15'h5760: q<=8'h4e;
	15'h5761: q<=8'h84;
	15'h5762: q<=8'h4f;
	15'h5763: q<=8'ha5;
	15'h5764: q<=8'hb4;
	15'h5765: q<=8'ha4;
	15'h5766: q<=8'h13;
	15'h5767: q<=8'h10;
	15'h5768: q<=8'h02;
	15'h5769: q<=8'h09;
	15'h576a: q<=8'h04;
	15'h576b: q<=8'ha4;
	15'h576c: q<=8'h14;
	15'h576d: q<=8'h10;
	15'h576e: q<=8'h02;
	15'h576f: q<=8'h09;
	15'h5770: q<=8'h02;
	15'h5771: q<=8'ha4;
	15'h5772: q<=8'h15;
	15'h5773: q<=8'h10;
	15'h5774: q<=8'h02;
	15'h5775: q<=8'h09;
	15'h5776: q<=8'h01;
	15'h5777: q<=8'h8d;
	15'h5778: q<=8'h00;
	15'h5779: q<=8'h40;
	15'h577a: q<=8'ha6;
	15'h577b: q<=8'h3e;
	15'h577c: q<=8'he8;
	15'h577d: q<=8'ha4;
	15'h577e: q<=8'h05;
	15'h577f: q<=8'hd0;
	15'h5780: q<=8'h10;
	15'h5781: q<=8'ha2;
	15'h5782: q<=8'h00;
	15'h5783: q<=8'ha4;
	15'h5784: q<=8'h07;
	15'h5785: q<=8'hc0;
	15'h5786: q<=8'h40;
	15'h5787: q<=8'h90;
	15'h5788: q<=8'h08;
	15'h5789: q<=8'ha6;
	15'h578a: q<=8'h06;
	15'h578b: q<=8'he0;
	15'h578c: q<=8'h02;
	15'h578d: q<=8'h90;
	15'h578e: q<=8'h02;
	15'h578f: q<=8'ha2;
	15'h5790: q<=8'h03;
	15'h5791: q<=8'hbd;
	15'h5792: q<=8'hdd;
	15'h5793: q<=8'hd7;
	15'h5794: q<=8'h45;
	15'h5795: q<=8'ha1;
	15'h5796: q<=8'h29;
	15'h5797: q<=8'h03;
	15'h5798: q<=8'h45;
	15'h5799: q<=8'ha1;
	15'h579a: q<=8'h85;
	15'h579b: q<=8'ha1;
	15'h579c: q<=8'h8d;
	15'h579d: q<=8'he0;
	15'h579e: q<=8'h60;
	15'h579f: q<=8'h20;
	15'h57a0: q<=8'h24;
	15'h57a1: q<=8'hcf;
	15'h57a2: q<=8'h20;
	15'h57a3: q<=8'h0a;
	15'h57a4: q<=8'hcd;
	15'h57a5: q<=8'he6;
	15'h57a6: q<=8'h53;
	15'h57a7: q<=8'he6;
	15'h57a8: q<=8'h07;
	15'h57a9: q<=8'hd0;
	15'h57aa: q<=8'h1e;
	15'h57ab: q<=8'hee;
	15'h57ac: q<=8'h06;
	15'h57ad: q<=8'h04;
	15'h57ae: q<=8'hd0;
	15'h57af: q<=8'h08;
	15'h57b0: q<=8'hee;
	15'h57b1: q<=8'h07;
	15'h57b2: q<=8'h04;
	15'h57b3: q<=8'hd0;
	15'h57b4: q<=8'h03;
	15'h57b5: q<=8'hee;
	15'h57b6: q<=8'h08;
	15'h57b7: q<=8'h04;
	15'h57b8: q<=8'h24;
	15'h57b9: q<=8'h05;
	15'h57ba: q<=8'h50;
	15'h57bb: q<=8'h0d;
	15'h57bc: q<=8'hee;
	15'h57bd: q<=8'h09;
	15'h57be: q<=8'h04;
	15'h57bf: q<=8'hd0;
	15'h57c0: q<=8'h08;
	15'h57c1: q<=8'hee;
	15'h57c2: q<=8'h0a;
	15'h57c3: q<=8'h04;
	15'h57c4: q<=8'hd0;
	15'h57c5: q<=8'h03;
	15'h57c6: q<=8'hee;
	15'h57c7: q<=8'h0b;
	15'h57c8: q<=8'h04;
	15'h57c9: q<=8'h2c;
	15'h57ca: q<=8'h00;
	15'h57cb: q<=8'h0c;
	15'h57cc: q<=8'h50;
	15'h57cd: q<=8'h09;
	15'h57ce: q<=8'hee;
	15'h57cf: q<=8'h33;
	15'h57d0: q<=8'h01;
	15'h57d1: q<=8'h8d;
	15'h57d2: q<=8'h00;
	15'h57d3: q<=8'h58;
	15'h57d4: q<=8'h8d;
	15'h57d5: q<=8'h00;
	15'h57d6: q<=8'h48;
	15'h57d7: q<=8'h68;
	15'h57d8: q<=8'ha8;
	15'h57d9: q<=8'h68;
	15'h57da: q<=8'haa;
	15'h57db: q<=8'h68;
	15'h57dc: q<=8'h40;
	15'h57dd: q<=8'hff;
	15'h57de: q<=8'hfd;
	15'h57df: q<=8'hfe;
	15'h57e0: q<=8'hfc;
	15'h57e1: q<=8'ha9;
	15'h57e2: q<=8'h00;
	15'h57e3: q<=8'h85;
	15'h57e4: q<=8'h05;
	15'h57e5: q<=8'ha9;
	15'h57e6: q<=8'h02;
	15'h57e7: q<=8'h85;
	15'h57e8: q<=8'h01;
	15'h57e9: q<=8'had;
	15'h57ea: q<=8'hca;
	15'h57eb: q<=8'h01;
	15'h57ec: q<=8'hd0;
	15'h57ed: q<=8'h15;
	15'h57ee: q<=8'had;
	15'h57ef: q<=8'h00;
	15'h57f0: q<=8'h0c;
	15'h57f1: q<=8'h29;
	15'h57f2: q<=8'h10;
	15'h57f3: q<=8'hf0;
	15'h57f4: q<=8'h0e;
	15'h57f5: q<=8'ha9;
	15'h57f6: q<=8'h00;
	15'h57f7: q<=8'h85;
	15'h57f8: q<=8'h00;
	15'h57f9: q<=8'had;
	15'h57fa: q<=8'hc9;
	15'h57fb: q<=8'h01;
	15'h57fc: q<=8'h29;
	15'h57fd: q<=8'h03;
	15'h57fe: q<=8'hf0;
	15'h57ff: q<=8'h03;
	15'h5800: q<=8'h20;
	15'h5801: q<=8'hac;
	15'h5802: q<=8'hab;
	15'h5803: q<=8'h60;
	15'h5804: q<=8'h20;
	15'h5805: q<=8'hbb;
	15'h5806: q<=8'hd6;
	15'h5807: q<=8'h20;
	15'h5808: q<=8'ha8;
	15'h5809: q<=8'haa;
	15'h580a: q<=8'h20;
	15'h580b: q<=8'h0d;
	15'h580c: q<=8'hdd;
	15'h580d: q<=8'h20;
	15'h580e: q<=8'h41;
	15'h580f: q<=8'hdd;
	15'h5810: q<=8'had;
	15'h5811: q<=8'h58;
	15'h5812: q<=8'h01;
	15'h5813: q<=8'h85;
	15'h5814: q<=8'h37;
	15'h5815: q<=8'h20;
	15'h5816: q<=8'h53;
	15'h5817: q<=8'hdf;
	15'h5818: q<=8'ha9;
	15'h5819: q<=8'he8;
	15'h581a: q<=8'ha2;
	15'h581b: q<=8'hc0;
	15'h581c: q<=8'h20;
	15'h581d: q<=8'h75;
	15'h581e: q<=8'hdf;
	15'h581f: q<=8'ha9;
	15'h5820: q<=8'h32;
	15'h5821: q<=8'ha2;
	15'h5822: q<=8'h6c;
	15'h5823: q<=8'h20;
	15'h5824: q<=8'h39;
	15'h5825: q<=8'hdf;
	15'h5826: q<=8'hc6;
	15'h5827: q<=8'h37;
	15'h5828: q<=8'hd0;
	15'h5829: q<=8'hf5;
	15'h582a: q<=8'had;
	15'h582b: q<=8'h6a;
	15'h582c: q<=8'h01;
	15'h582d: q<=8'h29;
	15'h582e: q<=8'h03;
	15'h582f: q<=8'h0a;
	15'h5830: q<=8'ha8;
	15'h5831: q<=8'hb9;
	15'h5832: q<=8'h1f;
	15'h5833: q<=8'h3f;
	15'h5834: q<=8'hbe;
	15'h5835: q<=8'h1e;
	15'h5836: q<=8'h3f;
	15'h5837: q<=8'h20;
	15'h5838: q<=8'h39;
	15'h5839: q<=8'hdf;
	15'h583a: q<=8'had;
	15'h583b: q<=8'h00;
	15'h583c: q<=8'h02;
	15'h583d: q<=8'h20;
	15'h583e: q<=8'hce;
	15'h583f: q<=8'had;
	15'h5840: q<=8'h8d;
	15'h5841: q<=8'h00;
	15'h5842: q<=8'h02;
	15'h5843: q<=8'h29;
	15'h5844: q<=8'h06;
	15'h5845: q<=8'h48;
	15'h5846: q<=8'ha8;
	15'h5847: q<=8'hb9;
	15'h5848: q<=8'h17;
	15'h5849: q<=8'h3f;
	15'h584a: q<=8'hbe;
	15'h584b: q<=8'h16;
	15'h584c: q<=8'h3f;
	15'h584d: q<=8'h20;
	15'h584e: q<=8'h39;
	15'h584f: q<=8'hdf;
	15'h5850: q<=8'h68;
	15'h5851: q<=8'h4a;
	15'h5852: q<=8'haa;
	15'h5853: q<=8'ha5;
	15'h5854: q<=8'h4d;
	15'h5855: q<=8'h3d;
	15'h5856: q<=8'hb6;
	15'h5857: q<=8'hd8;
	15'h5858: q<=8'hdd;
	15'h5859: q<=8'hb6;
	15'h585a: q<=8'hd8;
	15'h585b: q<=8'hd0;
	15'h585c: q<=8'h1a;
	15'h585d: q<=8'hca;
	15'h585e: q<=8'hca;
	15'h585f: q<=8'h10;
	15'h5860: q<=8'h03;
	15'h5861: q<=8'h4c;
	15'h5862: q<=8'h3f;
	15'h5863: q<=8'hd9;
	15'h5864: q<=8'hd0;
	15'h5865: q<=8'h06;
	15'h5866: q<=8'h20;
	15'h5867: q<=8'he9;
	15'h5868: q<=8'hdd;
	15'h5869: q<=8'hb8;
	15'h586a: q<=8'h50;
	15'h586b: q<=8'h0b;
	15'h586c: q<=8'h20;
	15'h586d: q<=8'hed;
	15'h586e: q<=8'hdd;
	15'h586f: q<=8'had;
	15'h5870: q<=8'hc9;
	15'h5871: q<=8'h01;
	15'h5872: q<=8'h09;
	15'h5873: q<=8'h03;
	15'h5874: q<=8'h8d;
	15'h5875: q<=8'hc9;
	15'h5876: q<=8'h01;
	15'h5877: q<=8'had;
	15'h5878: q<=8'hca;
	15'h5879: q<=8'h01;
	15'h587a: q<=8'h2d;
	15'h587b: q<=8'hc6;
	15'h587c: q<=8'h01;
	15'h587d: q<=8'hf0;
	15'h587e: q<=8'h07;
	15'h587f: q<=8'ha9;
	15'h5880: q<=8'h34;
	15'h5881: q<=8'ha2;
	15'h5882: q<=8'h6e;
	15'h5883: q<=8'h20;
	15'h5884: q<=8'h39;
	15'h5885: q<=8'hdf;
	15'h5886: q<=8'h20;
	15'h5887: q<=8'h53;
	15'h5888: q<=8'hdf;
	15'h5889: q<=8'ha5;
	15'h588a: q<=8'h09;
	15'h588b: q<=8'h29;
	15'h588c: q<=8'h1c;
	15'h588d: q<=8'h4a;
	15'h588e: q<=8'h4a;
	15'h588f: q<=8'haa;
	15'h5890: q<=8'hbd;
	15'h5891: q<=8'hba;
	15'h5892: q<=8'hd8;
	15'h5893: q<=8'ha0;
	15'h5894: q<=8'hee;
	15'h5895: q<=8'ha2;
	15'h5896: q<=8'h1b;
	15'h5897: q<=8'h20;
	15'h5898: q<=8'ha9;
	15'h5899: q<=8'hd8;
	15'h589a: q<=8'ha5;
	15'h589b: q<=8'h09;
	15'h589c: q<=8'h4a;
	15'h589d: q<=8'h4a;
	15'h589e: q<=8'h4a;
	15'h589f: q<=8'h4a;
	15'h58a0: q<=8'h4a;
	15'h58a1: q<=8'haa;
	15'h58a2: q<=8'hbd;
	15'h58a3: q<=8'hc2;
	15'h58a4: q<=8'hd8;
	15'h58a5: q<=8'ha0;
	15'h58a6: q<=8'h32;
	15'h58a7: q<=8'ha2;
	15'h58a8: q<=8'hf8;
	15'h58a9: q<=8'h85;
	15'h58aa: q<=8'h29;
	15'h58ab: q<=8'h98;
	15'h58ac: q<=8'h20;
	15'h58ad: q<=8'h75;
	15'h58ae: q<=8'hdf;
	15'h58af: q<=8'ha9;
	15'h58b0: q<=8'h29;
	15'h58b1: q<=8'ha0;
	15'h58b2: q<=8'h01;
	15'h58b3: q<=8'h4c;
	15'h58b4: q<=8'hb1;
	15'h58b5: q<=8'hdf;
	15'h58b6: q<=8'h18;
	15'h58b7: q<=8'h18;
	15'h58b8: q<=8'h30;
	15'h58b9: q<=8'h50;
	15'h58ba: q<=8'h11;
	15'h58bb: q<=8'h14;
	15'h58bc: q<=8'h15;
	15'h58bd: q<=8'h16;
	15'h58be: q<=8'h21;
	15'h58bf: q<=8'h24;
	15'h58c0: q<=8'h25;
	15'h58c1: q<=8'h26;
	15'h58c2: q<=8'h00;
	15'h58c3: q<=8'h12;
	15'h58c4: q<=8'h14;
	15'h58c5: q<=8'h24;
	15'h58c6: q<=8'h15;
	15'h58c7: q<=8'h13;
	15'h58c8: q<=8'h00;
	15'h58c9: q<=8'h00;
	15'h58ca: q<=8'ha8;
	15'h58cb: q<=8'ha9;
	15'h58cc: q<=8'h00;
	15'h58cd: q<=8'h84;
	15'h58ce: q<=8'h79;
	15'h58cf: q<=8'h4a;
	15'h58d0: q<=8'h4a;
	15'h58d1: q<=8'h0a;
	15'h58d2: q<=8'haa;
	15'h58d3: q<=8'h98;
	15'h58d4: q<=8'h29;
	15'h58d5: q<=8'h0f;
	15'h58d6: q<=8'hd0;
	15'h58d7: q<=8'h01;
	15'h58d8: q<=8'he8;
	15'h58d9: q<=8'h9a;
	15'h58da: q<=8'ha9;
	15'h58db: q<=8'ha2;
	15'h58dc: q<=8'h8d;
	15'h58dd: q<=8'hc1;
	15'h58de: q<=8'h60;
	15'h58df: q<=8'hba;
	15'h58e0: q<=8'hd0;
	15'h58e1: q<=8'h07;
	15'h58e2: q<=8'ha9;
	15'h58e3: q<=8'h60;
	15'h58e4: q<=8'ha0;
	15'h58e5: q<=8'h09;
	15'h58e6: q<=8'hb8;
	15'h58e7: q<=8'h50;
	15'h58e8: q<=8'h04;
	15'h58e9: q<=8'ha9;
	15'h58ea: q<=8'hc0;
	15'h58eb: q<=8'ha0;
	15'h58ec: q<=8'h01;
	15'h58ed: q<=8'h8d;
	15'h58ee: q<=8'hc0;
	15'h58ef: q<=8'h60;
	15'h58f0: q<=8'ha9;
	15'h58f1: q<=8'h03;
	15'h58f2: q<=8'h8d;
	15'h58f3: q<=8'he0;
	15'h58f4: q<=8'h60;
	15'h58f5: q<=8'ha2;
	15'h58f6: q<=8'h00;
	15'h58f7: q<=8'h2c;
	15'h58f8: q<=8'h00;
	15'h58f9: q<=8'h0c;
	15'h58fa: q<=8'h30;
	15'h58fb: q<=8'hfb;
	15'h58fc: q<=8'h2c;
	15'h58fd: q<=8'h00;
	15'h58fe: q<=8'h0c;
	15'h58ff: q<=8'h10;
	15'h5900: q<=8'hfb;
	15'h5901: q<=8'h8d;
	15'h5902: q<=8'h00;
	15'h5903: q<=8'h50;
	15'h5904: q<=8'hca;
	15'h5905: q<=8'hd0;
	15'h5906: q<=8'hf0;
	15'h5907: q<=8'h88;
	15'h5908: q<=8'hd0;
	15'h5909: q<=8'hed;
	15'h590a: q<=8'h8e;
	15'h590b: q<=8'hc1;
	15'h590c: q<=8'h60;
	15'h590d: q<=8'ha9;
	15'h590e: q<=8'h00;
	15'h590f: q<=8'h8d;
	15'h5910: q<=8'he0;
	15'h5911: q<=8'h60;
	15'h5912: q<=8'ha0;
	15'h5913: q<=8'h09;
	15'h5914: q<=8'h2c;
	15'h5915: q<=8'h00;
	15'h5916: q<=8'h0c;
	15'h5917: q<=8'h30;
	15'h5918: q<=8'hfb;
	15'h5919: q<=8'h2c;
	15'h591a: q<=8'h00;
	15'h591b: q<=8'h0c;
	15'h591c: q<=8'h10;
	15'h591d: q<=8'hfb;
	15'h591e: q<=8'h8d;
	15'h591f: q<=8'h00;
	15'h5920: q<=8'h50;
	15'h5921: q<=8'hca;
	15'h5922: q<=8'hd0;
	15'h5923: q<=8'hf0;
	15'h5924: q<=8'h88;
	15'h5925: q<=8'hd0;
	15'h5926: q<=8'hed;
	15'h5927: q<=8'hba;
	15'h5928: q<=8'hca;
	15'h5929: q<=8'h9a;
	15'h592a: q<=8'h10;
	15'h592b: q<=8'hae;
	15'h592c: q<=8'h4c;
	15'h592d: q<=8'h0a;
	15'h592e: q<=8'hda;
	15'h592f: q<=8'h51;
	15'h5930: q<=8'h00;
	15'h5931: q<=8'ha8;
	15'h5932: q<=8'ha5;
	15'h5933: q<=8'h01;
	15'h5934: q<=8'hc9;
	15'h5935: q<=8'h20;
	15'h5936: q<=8'h90;
	15'h5937: q<=8'h02;
	15'h5938: q<=8'he9;
	15'h5939: q<=8'h18;
	15'h593a: q<=8'h29;
	15'h593b: q<=8'h1f;
	15'h593c: q<=8'h4c;
	15'h593d: q<=8'hcd;
	15'h593e: q<=8'hd8;
	15'h593f: q<=8'h78;
	15'h5940: q<=8'h8d;
	15'h5941: q<=8'h00;
	15'h5942: q<=8'h50;
	15'h5943: q<=8'h8d;
	15'h5944: q<=8'h00;
	15'h5945: q<=8'h58;
	15'h5946: q<=8'ha2;
	15'h5947: q<=8'hff;
	15'h5948: q<=8'h9a;
	15'h5949: q<=8'hd8;
	15'h594a: q<=8'he8;
	15'h594b: q<=8'h8a;
	15'h594c: q<=8'ha8;
	15'h594d: q<=8'h84;
	15'h594e: q<=8'h00;
	15'h594f: q<=8'h86;
	15'h5950: q<=8'h01;
	15'h5951: q<=8'ha0;
	15'h5952: q<=8'h00;
	15'h5953: q<=8'h91;
	15'h5954: q<=8'h00;
	15'h5955: q<=8'hc8;
	15'h5956: q<=8'hd0;
	15'h5957: q<=8'hfb;
	15'h5958: q<=8'he8;
	15'h5959: q<=8'he0;
	15'h595a: q<=8'h08;
	15'h595b: q<=8'hd0;
	15'h595c: q<=8'h02;
	15'h595d: q<=8'ha2;
	15'h595e: q<=8'h20;
	15'h595f: q<=8'he0;
	15'h5960: q<=8'h30;
	15'h5961: q<=8'h8d;
	15'h5962: q<=8'h00;
	15'h5963: q<=8'h50;
	15'h5964: q<=8'h90;
	15'h5965: q<=8'he7;
	15'h5966: q<=8'h85;
	15'h5967: q<=8'h01;
	15'h5968: q<=8'h8d;
	15'h5969: q<=8'he0;
	15'h596a: q<=8'h60;
	15'h596b: q<=8'h8d;
	15'h596c: q<=8'hcf;
	15'h596d: q<=8'h60;
	15'h596e: q<=8'h8d;
	15'h596f: q<=8'hdf;
	15'h5970: q<=8'h60;
	15'h5971: q<=8'ha2;
	15'h5972: q<=8'h07;
	15'h5973: q<=8'h8e;
	15'h5974: q<=8'hcf;
	15'h5975: q<=8'h60;
	15'h5976: q<=8'h8e;
	15'h5977: q<=8'hdf;
	15'h5978: q<=8'h60;
	15'h5979: q<=8'he8;
	15'h597a: q<=8'h9d;
	15'h597b: q<=8'hc0;
	15'h597c: q<=8'h60;
	15'h597d: q<=8'h9d;
	15'h597e: q<=8'hd0;
	15'h597f: q<=8'h60;
	15'h5980: q<=8'hca;
	15'h5981: q<=8'h10;
	15'h5982: q<=8'hf7;
	15'h5983: q<=8'had;
	15'h5984: q<=8'h00;
	15'h5985: q<=8'h0c;
	15'h5986: q<=8'h29;
	15'h5987: q<=8'h10;
	15'h5988: q<=8'hf0;
	15'h5989: q<=8'h1f;
	15'h598a: q<=8'h8d;
	15'h598b: q<=8'h00;
	15'h598c: q<=8'h50;
	15'h598d: q<=8'hce;
	15'h598e: q<=8'h00;
	15'h598f: q<=8'h01;
	15'h5990: q<=8'hd0;
	15'h5991: q<=8'hf8;
	15'h5992: q<=8'hce;
	15'h5993: q<=8'h01;
	15'h5994: q<=8'h01;
	15'h5995: q<=8'hd0;
	15'h5996: q<=8'hf3;
	15'h5997: q<=8'ha9;
	15'h5998: q<=8'h10;
	15'h5999: q<=8'h85;
	15'h599a: q<=8'hb4;
	15'h599b: q<=8'h20;
	15'h599c: q<=8'h11;
	15'h599d: q<=8'hde;
	15'h599e: q<=8'h20;
	15'h599f: q<=8'hac;
	15'h59a0: q<=8'hab;
	15'h59a1: q<=8'h20;
	15'h59a2: q<=8'h6e;
	15'h59a3: q<=8'hc1;
	15'h59a4: q<=8'h58;
	15'h59a5: q<=8'h4c;
	15'h59a6: q<=8'ha0;
	15'h59a7: q<=8'hc7;
	15'h59a8: q<=8'ha0;
	15'h59a9: q<=8'ha2;
	15'h59aa: q<=8'h11;
	15'h59ab: q<=8'h9a;
	15'h59ac: q<=8'ha0;
	15'h59ad: q<=8'h00;
	15'h59ae: q<=8'hba;
	15'h59af: q<=8'h96;
	15'h59b0: q<=8'h00;
	15'h59b1: q<=8'ha2;
	15'h59b2: q<=8'h01;
	15'h59b3: q<=8'hc8;
	15'h59b4: q<=8'hb9;
	15'h59b5: q<=8'h00;
	15'h59b6: q<=8'h00;
	15'h59b7: q<=8'hf0;
	15'h59b8: q<=8'h03;
	15'h59b9: q<=8'h4c;
	15'h59ba: q<=8'hca;
	15'h59bb: q<=8'hd8;
	15'h59bc: q<=8'he8;
	15'h59bd: q<=8'hd0;
	15'h59be: q<=8'hf4;
	15'h59bf: q<=8'hba;
	15'h59c0: q<=8'h8a;
	15'h59c1: q<=8'h8d;
	15'h59c2: q<=8'h00;
	15'h59c3: q<=8'h50;
	15'h59c4: q<=8'hc8;
	15'h59c5: q<=8'h59;
	15'h59c6: q<=8'h00;
	15'h59c7: q<=8'h00;
	15'h59c8: q<=8'hd0;
	15'h59c9: q<=8'hef;
	15'h59ca: q<=8'h99;
	15'h59cb: q<=8'h00;
	15'h59cc: q<=8'h00;
	15'h59cd: q<=8'hc8;
	15'h59ce: q<=8'hd0;
	15'h59cf: q<=8'hde;
	15'h59d0: q<=8'hba;
	15'h59d1: q<=8'h8a;
	15'h59d2: q<=8'h0a;
	15'h59d3: q<=8'haa;
	15'h59d4: q<=8'h90;
	15'h59d5: q<=8'hd5;
	15'h59d6: q<=8'ha0;
	15'h59d7: q<=8'h00;
	15'h59d8: q<=8'ha2;
	15'h59d9: q<=8'h01;
	15'h59da: q<=8'h84;
	15'h59db: q<=8'h00;
	15'h59dc: q<=8'h86;
	15'h59dd: q<=8'h01;
	15'h59de: q<=8'ha0;
	15'h59df: q<=8'h00;
	15'h59e0: q<=8'hb1;
	15'h59e1: q<=8'h00;
	15'h59e2: q<=8'hf0;
	15'h59e3: q<=8'h03;
	15'h59e4: q<=8'h4c;
	15'h59e5: q<=8'h31;
	15'h59e6: q<=8'hd9;
	15'h59e7: q<=8'ha9;
	15'h59e8: q<=8'h11;
	15'h59e9: q<=8'h91;
	15'h59ea: q<=8'h00;
	15'h59eb: q<=8'hd1;
	15'h59ec: q<=8'h00;
	15'h59ed: q<=8'hf0;
	15'h59ee: q<=8'h03;
	15'h59ef: q<=8'h4c;
	15'h59f0: q<=8'h2f;
	15'h59f1: q<=8'hd9;
	15'h59f2: q<=8'h0a;
	15'h59f3: q<=8'h90;
	15'h59f4: q<=8'hf4;
	15'h59f5: q<=8'ha9;
	15'h59f6: q<=8'h00;
	15'h59f7: q<=8'h91;
	15'h59f8: q<=8'h00;
	15'h59f9: q<=8'hc8;
	15'h59fa: q<=8'hd0;
	15'h59fb: q<=8'he4;
	15'h59fc: q<=8'h8d;
	15'h59fd: q<=8'h00;
	15'h59fe: q<=8'h50;
	15'h59ff: q<=8'he8;
	15'h5a00: q<=8'he0;
	15'h5a01: q<=8'h08;
	15'h5a02: q<=8'hd0;
	15'h5a03: q<=8'h02;
	15'h5a04: q<=8'ha2;
	15'h5a05: q<=8'h20;
	15'h5a06: q<=8'he0;
	15'h5a07: q<=8'h30;
	15'h5a08: q<=8'h90;
	15'h5a09: q<=8'hd0;
	15'h5a0a: q<=8'ha9;
	15'h5a0b: q<=8'h00;
	15'h5a0c: q<=8'ha8;
	15'h5a0d: q<=8'haa;
	15'h5a0e: q<=8'h85;
	15'h5a0f: q<=8'h3b;
	15'h5a10: q<=8'ha9;
	15'h5a11: q<=8'h30;
	15'h5a12: q<=8'h85;
	15'h5a13: q<=8'h3c;
	15'h5a14: q<=8'ha9;
	15'h5a15: q<=8'h08;
	15'h5a16: q<=8'h85;
	15'h5a17: q<=8'h38;
	15'h5a18: q<=8'h8a;
	15'h5a19: q<=8'h51;
	15'h5a1a: q<=8'h3b;
	15'h5a1b: q<=8'hc8;
	15'h5a1c: q<=8'hd0;
	15'h5a1d: q<=8'hfb;
	15'h5a1e: q<=8'he6;
	15'h5a1f: q<=8'h3c;
	15'h5a20: q<=8'h8d;
	15'h5a21: q<=8'h00;
	15'h5a22: q<=8'h50;
	15'h5a23: q<=8'hc6;
	15'h5a24: q<=8'h38;
	15'h5a25: q<=8'hd0;
	15'h5a26: q<=8'hf2;
	15'h5a27: q<=8'h95;
	15'h5a28: q<=8'h7d;
	15'h5a29: q<=8'he8;
	15'h5a2a: q<=8'he0;
	15'h5a2b: q<=8'h02;
	15'h5a2c: q<=8'hd0;
	15'h5a2d: q<=8'h04;
	15'h5a2e: q<=8'ha9;
	15'h5a2f: q<=8'h90;
	15'h5a30: q<=8'h85;
	15'h5a31: q<=8'h3c;
	15'h5a32: q<=8'he0;
	15'h5a33: q<=8'h0c;
	15'h5a34: q<=8'h90;
	15'h5a35: q<=8'hde;
	15'h5a36: q<=8'ha5;
	15'h5a37: q<=8'h7d;
	15'h5a38: q<=8'hf0;
	15'h5a39: q<=8'h0a;
	15'h5a3a: q<=8'ha9;
	15'h5a3b: q<=8'h40;
	15'h5a3c: q<=8'ha2;
	15'h5a3d: q<=8'ha4;
	15'h5a3e: q<=8'h8d;
	15'h5a3f: q<=8'hc4;
	15'h5a40: q<=8'h60;
	15'h5a41: q<=8'h8e;
	15'h5a42: q<=8'hc5;
	15'h5a43: q<=8'h60;
	15'h5a44: q<=8'ha2;
	15'h5a45: q<=8'h05;
	15'h5a46: q<=8'had;
	15'h5a47: q<=8'hca;
	15'h5a48: q<=8'h60;
	15'h5a49: q<=8'hcd;
	15'h5a4a: q<=8'hca;
	15'h5a4b: q<=8'h60;
	15'h5a4c: q<=8'hd0;
	15'h5a4d: q<=8'h05;
	15'h5a4e: q<=8'hca;
	15'h5a4f: q<=8'h10;
	15'h5a50: q<=8'hf8;
	15'h5a51: q<=8'h85;
	15'h5a52: q<=8'h7a;
	15'h5a53: q<=8'ha2;
	15'h5a54: q<=8'h05;
	15'h5a55: q<=8'had;
	15'h5a56: q<=8'hda;
	15'h5a57: q<=8'h60;
	15'h5a58: q<=8'hcd;
	15'h5a59: q<=8'hda;
	15'h5a5a: q<=8'h60;
	15'h5a5b: q<=8'hd0;
	15'h5a5c: q<=8'h05;
	15'h5a5d: q<=8'hca;
	15'h5a5e: q<=8'h10;
	15'h5a5f: q<=8'hf8;
	15'h5a60: q<=8'h85;
	15'h5a61: q<=8'h7b;
	15'h5a62: q<=8'h20;
	15'h5a63: q<=8'h11;
	15'h5a64: q<=8'hde;
	15'h5a65: q<=8'ha0;
	15'h5a66: q<=8'h02;
	15'h5a67: q<=8'had;
	15'h5a68: q<=8'hc9;
	15'h5a69: q<=8'h01;
	15'h5a6a: q<=8'hf0;
	15'h5a6b: q<=8'h0a;
	15'h5a6c: q<=8'h85;
	15'h5a6d: q<=8'h7c;
	15'h5a6e: q<=8'h20;
	15'h5a6f: q<=8'hf1;
	15'h5a70: q<=8'hdd;
	15'h5a71: q<=8'ha0;
	15'h5a72: q<=8'h00;
	15'h5a73: q<=8'h8c;
	15'h5a74: q<=8'hc9;
	15'h5a75: q<=8'h01;
	15'h5a76: q<=8'h84;
	15'h5a77: q<=8'h00;
	15'h5a78: q<=8'ha2;
	15'h5a79: q<=8'h07;
	15'h5a7a: q<=8'hbd;
	15'h5a7b: q<=8'hf9;
	15'h5a7c: q<=8'hda;
	15'h5a7d: q<=8'h9d;
	15'h5a7e: q<=8'h00;
	15'h5a7f: q<=8'h08;
	15'h5a80: q<=8'hca;
	15'h5a81: q<=8'h10;
	15'h5a82: q<=8'hf7;
	15'h5a83: q<=8'ha9;
	15'h5a84: q<=8'h00;
	15'h5a85: q<=8'h8d;
	15'h5a86: q<=8'he0;
	15'h5a87: q<=8'h60;
	15'h5a88: q<=8'ha9;
	15'h5a89: q<=8'h10;
	15'h5a8a: q<=8'h8d;
	15'h5a8b: q<=8'h00;
	15'h5a8c: q<=8'h40;
	15'h5a8d: q<=8'ha0;
	15'h5a8e: q<=8'h04;
	15'h5a8f: q<=8'ha2;
	15'h5a90: q<=8'h14;
	15'h5a91: q<=8'h2c;
	15'h5a92: q<=8'h00;
	15'h5a93: q<=8'h0c;
	15'h5a94: q<=8'h10;
	15'h5a95: q<=8'hfb;
	15'h5a96: q<=8'h2c;
	15'h5a97: q<=8'h00;
	15'h5a98: q<=8'h0c;
	15'h5a99: q<=8'h30;
	15'h5a9a: q<=8'hfb;
	15'h5a9b: q<=8'hca;
	15'h5a9c: q<=8'h10;
	15'h5a9d: q<=8'hf3;
	15'h5a9e: q<=8'h88;
	15'h5a9f: q<=8'h30;
	15'h5aa0: q<=8'h08;
	15'h5aa1: q<=8'h8d;
	15'h5aa2: q<=8'h00;
	15'h5aa3: q<=8'h50;
	15'h5aa4: q<=8'h2c;
	15'h5aa5: q<=8'h00;
	15'h5aa6: q<=8'h0c;
	15'h5aa7: q<=8'h50;
	15'h5aa8: q<=8'he6;
	15'h5aa9: q<=8'h8d;
	15'h5aaa: q<=8'h00;
	15'h5aab: q<=8'h58;
	15'h5aac: q<=8'ha9;
	15'h5aad: q<=8'h00;
	15'h5aae: q<=8'h85;
	15'h5aaf: q<=8'h74;
	15'h5ab0: q<=8'ha9;
	15'h5ab1: q<=8'h20;
	15'h5ab2: q<=8'h85;
	15'h5ab3: q<=8'h75;
	15'h5ab4: q<=8'h8d;
	15'h5ab5: q<=8'hcb;
	15'h5ab6: q<=8'h60;
	15'h5ab7: q<=8'had;
	15'h5ab8: q<=8'hc8;
	15'h5ab9: q<=8'h60;
	15'h5aba: q<=8'h85;
	15'h5abb: q<=8'h52;
	15'h5abc: q<=8'h29;
	15'h5abd: q<=8'h0f;
	15'h5abe: q<=8'h85;
	15'h5abf: q<=8'h50;
	15'h5ac0: q<=8'had;
	15'h5ac1: q<=8'h00;
	15'h5ac2: q<=8'h0c;
	15'h5ac3: q<=8'h49;
	15'h5ac4: q<=8'hff;
	15'h5ac5: q<=8'h29;
	15'h5ac6: q<=8'h2f;
	15'h5ac7: q<=8'h85;
	15'h5ac8: q<=8'h4e;
	15'h5ac9: q<=8'h29;
	15'h5aca: q<=8'h28;
	15'h5acb: q<=8'hf0;
	15'h5acc: q<=8'h0b;
	15'h5acd: q<=8'h06;
	15'h5ace: q<=8'h4c;
	15'h5acf: q<=8'h90;
	15'h5ad0: q<=8'h04;
	15'h5ad1: q<=8'he6;
	15'h5ad2: q<=8'h00;
	15'h5ad3: q<=8'he6;
	15'h5ad4: q<=8'h00;
	15'h5ad5: q<=8'hb8;
	15'h5ad6: q<=8'h50;
	15'h5ad7: q<=8'h04;
	15'h5ad8: q<=8'ha9;
	15'h5ad9: q<=8'h20;
	15'h5ada: q<=8'h85;
	15'h5adb: q<=8'h4c;
	15'h5adc: q<=8'h20;
	15'h5add: q<=8'h0f;
	15'h5ade: q<=8'hdb;
	15'h5adf: q<=8'h20;
	15'h5ae0: q<=8'h0d;
	15'h5ae1: q<=8'hdf;
	15'h5ae2: q<=8'h8d;
	15'h5ae3: q<=8'h00;
	15'h5ae4: q<=8'h48;
	15'h5ae5: q<=8'he6;
	15'h5ae6: q<=8'h03;
	15'h5ae7: q<=8'ha5;
	15'h5ae8: q<=8'h03;
	15'h5ae9: q<=8'h29;
	15'h5aea: q<=8'h03;
	15'h5aeb: q<=8'hd0;
	15'h5aec: q<=8'h03;
	15'h5aed: q<=8'h20;
	15'h5aee: q<=8'h1b;
	15'h5aef: q<=8'hde;
	15'h5af0: q<=8'had;
	15'h5af1: q<=8'h00;
	15'h5af2: q<=8'h0c;
	15'h5af3: q<=8'h29;
	15'h5af4: q<=8'h10;
	15'h5af5: q<=8'hf0;
	15'h5af6: q<=8'h96;
	15'h5af7: q<=8'hd0;
	15'h5af8: q<=8'hfe;
	15'h5af9: q<=8'h00;
	15'h5afa: q<=8'h04;
	15'h5afb: q<=8'h08;
	15'h5afc: q<=8'h0c;
	15'h5afd: q<=8'h03;
	15'h5afe: q<=8'h07;
	15'h5aff: q<=8'h0b;
	15'h5b00: q<=8'h0b;
	15'h5b01: q<=8'h59;
	15'h5b02: q<=8'hdb;
	15'h5b03: q<=8'hf6;
	15'h5b04: q<=8'hdb;
	15'h5b05: q<=8'h83;
	15'h5b06: q<=8'hdb;
	15'h5b07: q<=8'h99;
	15'h5b08: q<=8'hdb;
	15'h5b09: q<=8'h7d;
	15'h5b0a: q<=8'hdb;
	15'h5b0b: q<=8'h6e;
	15'h5b0c: q<=8'hdb;
	15'h5b0d: q<=8'h21;
	15'h5b0e: q<=8'hdb;
	15'h5b0f: q<=8'ha6;
	15'h5b10: q<=8'h00;
	15'h5b11: q<=8'he0;
	15'h5b12: q<=8'h0e;
	15'h5b13: q<=8'h90;
	15'h5b14: q<=8'h04;
	15'h5b15: q<=8'ha2;
	15'h5b16: q<=8'h02;
	15'h5b17: q<=8'h86;
	15'h5b18: q<=8'h00;
	15'h5b19: q<=8'hbd;
	15'h5b1a: q<=8'h02;
	15'h5b1b: q<=8'hdb;
	15'h5b1c: q<=8'h48;
	15'h5b1d: q<=8'hbd;
	15'h5b1e: q<=8'h01;
	15'h5b1f: q<=8'hdb;
	15'h5b20: q<=8'h48;
	15'h5b21: q<=8'h60;
	15'h5b22: q<=8'ha9;
	15'h5b23: q<=8'h00;
	15'h5b24: q<=8'h8d;
	15'h5b25: q<=8'he0;
	15'h5b26: q<=8'h60;
	15'h5b27: q<=8'h8d;
	15'h5b28: q<=8'h80;
	15'h5b29: q<=8'h60;
	15'h5b2a: q<=8'h8d;
	15'h5b2b: q<=8'hc0;
	15'h5b2c: q<=8'h60;
	15'h5b2d: q<=8'h8d;
	15'h5b2e: q<=8'hd0;
	15'h5b2f: q<=8'h60;
	15'h5b30: q<=8'h8d;
	15'h5b31: q<=8'h00;
	15'h5b32: q<=8'h60;
	15'h5b33: q<=8'h8d;
	15'h5b34: q<=8'h40;
	15'h5b35: q<=8'h60;
	15'h5b36: q<=8'had;
	15'h5b37: q<=8'h40;
	15'h5b38: q<=8'h60;
	15'h5b39: q<=8'had;
	15'h5b3a: q<=8'h60;
	15'h5b3b: q<=8'h60;
	15'h5b3c: q<=8'had;
	15'h5b3d: q<=8'h70;
	15'h5b3e: q<=8'h60;
	15'h5b3f: q<=8'had;
	15'h5b40: q<=8'h50;
	15'h5b41: q<=8'h60;
	15'h5b42: q<=8'ha9;
	15'h5b43: q<=8'h08;
	15'h5b44: q<=8'h8d;
	15'h5b45: q<=8'he0;
	15'h5b46: q<=8'h60;
	15'h5b47: q<=8'ha9;
	15'h5b48: q<=8'h01;
	15'h5b49: q<=8'ha2;
	15'h5b4a: q<=8'h1f;
	15'h5b4b: q<=8'h18;
	15'h5b4c: q<=8'h9d;
	15'h5b4d: q<=8'h80;
	15'h5b4e: q<=8'h60;
	15'h5b4f: q<=8'h2a;
	15'h5b50: q<=8'hca;
	15'h5b51: q<=8'h10;
	15'h5b52: q<=8'hf9;
	15'h5b53: q<=8'ha9;
	15'h5b54: q<=8'h34;
	15'h5b55: q<=8'ha2;
	15'h5b56: q<=8'ha6;
	15'h5b57: q<=8'h4c;
	15'h5b58: q<=8'h39;
	15'h5b59: q<=8'hdf;
	15'h5b5a: q<=8'had;
	15'h5b5b: q<=8'hca;
	15'h5b5c: q<=8'h01;
	15'h5b5d: q<=8'h0d;
	15'h5b5e: q<=8'hc7;
	15'h5b5f: q<=8'h01;
	15'h5b60: q<=8'hd0;
	15'h5b61: q<=8'h0c;
	15'h5b62: q<=8'h20;
	15'h5b63: q<=8'h11;
	15'h5b64: q<=8'hde;
	15'h5b65: q<=8'had;
	15'h5b66: q<=8'hc9;
	15'h5b67: q<=8'h01;
	15'h5b68: q<=8'h85;
	15'h5b69: q<=8'h7c;
	15'h5b6a: q<=8'ha9;
	15'h5b6b: q<=8'h02;
	15'h5b6c: q<=8'h85;
	15'h5b6d: q<=8'h00;
	15'h5b6e: q<=8'h60;
	15'h5b6f: q<=8'ha5;
	15'h5b70: q<=8'h50;
	15'h5b71: q<=8'h4a;
	15'h5b72: q<=8'ha8;
	15'h5b73: q<=8'ha9;
	15'h5b74: q<=8'h68;
	15'h5b75: q<=8'h20;
	15'h5b76: q<=8'h4c;
	15'h5b77: q<=8'hdf;
	15'h5b78: q<=8'ha2;
	15'h5b79: q<=8'h4e;
	15'h5b7a: q<=8'ha9;
	15'h5b7b: q<=8'h33;
	15'h5b7c: q<=8'hd0;
	15'h5b7d: q<=8'h0a;
	15'h5b7e: q<=8'ha2;
	15'h5b7f: q<=8'hb6;
	15'h5b80: q<=8'ha9;
	15'h5b81: q<=8'h32;
	15'h5b82: q<=8'hd0;
	15'h5b83: q<=8'h04;
	15'h5b84: q<=8'ha9;
	15'h5b85: q<=8'h33;
	15'h5b86: q<=8'ha2;
	15'h5b87: q<=8'h0a;
	15'h5b88: q<=8'h20;
	15'h5b89: q<=8'h39;
	15'h5b8a: q<=8'hdf;
	15'h5b8b: q<=8'ha2;
	15'h5b8c: q<=8'h06;
	15'h5b8d: q<=8'ha9;
	15'h5b8e: q<=8'h00;
	15'h5b8f: q<=8'h9d;
	15'h5b90: q<=8'hc1;
	15'h5b91: q<=8'h60;
	15'h5b92: q<=8'h9d;
	15'h5b93: q<=8'hd1;
	15'h5b94: q<=8'h60;
	15'h5b95: q<=8'hca;
	15'h5b96: q<=8'hca;
	15'h5b97: q<=8'h10;
	15'h5b98: q<=8'hf6;
	15'h5b99: q<=8'h60;
	15'h5b9a: q<=8'ha5;
	15'h5b9b: q<=8'h03;
	15'h5b9c: q<=8'h29;
	15'h5b9d: q<=8'h3f;
	15'h5b9e: q<=8'hd0;
	15'h5b9f: q<=8'h02;
	15'h5ba0: q<=8'he6;
	15'h5ba1: q<=8'h39;
	15'h5ba2: q<=8'ha5;
	15'h5ba3: q<=8'h39;
	15'h5ba4: q<=8'h29;
	15'h5ba5: q<=8'h07;
	15'h5ba6: q<=8'haa;
	15'h5ba7: q<=8'hbc;
	15'h5ba8: q<=8'hd5;
	15'h5ba9: q<=8'hdb;
	15'h5baa: q<=8'ha9;
	15'h5bab: q<=8'h00;
	15'h5bac: q<=8'h99;
	15'h5bad: q<=8'hc1;
	15'h5bae: q<=8'h60;
	15'h5baf: q<=8'hbc;
	15'h5bb0: q<=8'hd6;
	15'h5bb1: q<=8'hdb;
	15'h5bb2: q<=8'hbd;
	15'h5bb3: q<=8'hdc;
	15'h5bb4: q<=8'hdf;
	15'h5bb5: q<=8'h99;
	15'h5bb6: q<=8'hc0;
	15'h5bb7: q<=8'h60;
	15'h5bb8: q<=8'ha9;
	15'h5bb9: q<=8'ha8;
	15'h5bba: q<=8'h99;
	15'h5bbb: q<=8'hc1;
	15'h5bbc: q<=8'h60;
	15'h5bbd: q<=8'ha9;
	15'h5bbe: q<=8'h34;
	15'h5bbf: q<=8'ha2;
	15'h5bc0: q<=8'h56;
	15'h5bc1: q<=8'h20;
	15'h5bc2: q<=8'h39;
	15'h5bc3: q<=8'hdf;
	15'h5bc4: q<=8'ha5;
	15'h5bc5: q<=8'h03;
	15'h5bc6: q<=8'h29;
	15'h5bc7: q<=8'h7f;
	15'h5bc8: q<=8'ha8;
	15'h5bc9: q<=8'ha9;
	15'h5bca: q<=8'h01;
	15'h5bcb: q<=8'h20;
	15'h5bcc: q<=8'h6c;
	15'h5bcd: q<=8'hdf;
	15'h5bce: q<=8'ha9;
	15'h5bcf: q<=8'h34;
	15'h5bd0: q<=8'ha2;
	15'h5bd1: q<=8'haa;
	15'h5bd2: q<=8'h4c;
	15'h5bd3: q<=8'h39;
	15'h5bd4: q<=8'hdf;
	15'h5bd5: q<=8'h16;
	15'h5bd6: q<=8'h00;
	15'h5bd7: q<=8'h10;
	15'h5bd8: q<=8'h02;
	15'h5bd9: q<=8'h12;
	15'h5bda: q<=8'h04;
	15'h5bdb: q<=8'h14;
	15'h5bdc: q<=8'h06;
	15'h5bdd: q<=8'h16;
	15'h5bde: q<=8'h00;
	15'h5bdf: q<=8'hea;
	15'h5be0: q<=8'h8d;
	15'h5be1: q<=8'hdb;
	15'h5be2: q<=8'h60;
	15'h5be3: q<=8'had;
	15'h5be4: q<=8'hd8;
	15'h5be5: q<=8'h60;
	15'h5be6: q<=8'h29;
	15'h5be7: q<=8'h07;
	15'h5be8: q<=8'h85;
	15'h5be9: q<=8'h37;
	15'h5bea: q<=8'h8d;
	15'h5beb: q<=8'hcb;
	15'h5bec: q<=8'h60;
	15'h5bed: q<=8'had;
	15'h5bee: q<=8'hc8;
	15'h5bef: q<=8'h60;
	15'h5bf0: q<=8'h29;
	15'h5bf1: q<=8'h20;
	15'h5bf2: q<=8'h4a;
	15'h5bf3: q<=8'h4a;
	15'h5bf4: q<=8'h05;
	15'h5bf5: q<=8'h37;
	15'h5bf6: q<=8'h60;
	15'h5bf7: q<=8'ha5;
	15'h5bf8: q<=8'h2e;
	15'h5bf9: q<=8'hf0;
	15'h5bfa: q<=8'h1e;
	15'h5bfb: q<=8'h8d;
	15'h5bfc: q<=8'h95;
	15'h5bfd: q<=8'h60;
	15'h5bfe: q<=8'h8d;
	15'h5bff: q<=8'h8d;
	15'h5c00: q<=8'h60;
	15'h5c01: q<=8'ha5;
	15'h5c02: q<=8'h2f;
	15'h5c03: q<=8'h8d;
	15'h5c04: q<=8'h96;
	15'h5c05: q<=8'h60;
	15'h5c06: q<=8'ha2;
	15'h5c07: q<=8'h00;
	15'h5c08: q<=8'h20;
	15'h5c09: q<=8'he6;
	15'h5c0a: q<=8'hdc;
	15'h5c0b: q<=8'hc9;
	15'h5c0c: q<=8'h01;
	15'h5c0d: q<=8'hd0;
	15'h5c0e: q<=8'h06;
	15'h5c0f: q<=8'h98;
	15'h5c10: q<=8'hd0;
	15'h5c11: q<=8'h03;
	15'h5c12: q<=8'h8a;
	15'h5c13: q<=8'h10;
	15'h5c14: q<=8'h04;
	15'h5c15: q<=8'ha9;
	15'h5c16: q<=8'hff;
	15'h5c17: q<=8'h85;
	15'h5c18: q<=8'h78;
	15'h5c19: q<=8'ha2;
	15'h5c1a: q<=8'h00;
	15'h5c1b: q<=8'h86;
	15'h5c1c: q<=8'h73;
	15'h5c1d: q<=8'he6;
	15'h5c1e: q<=8'h2e;
	15'h5c1f: q<=8'hd0;
	15'h5c20: q<=8'h06;
	15'h5c21: q<=8'he6;
	15'h5c22: q<=8'h2f;
	15'h5c23: q<=8'h10;
	15'h5c24: q<=8'h02;
	15'h5c25: q<=8'h86;
	15'h5c26: q<=8'h2f;
	15'h5c27: q<=8'h8d;
	15'h5c28: q<=8'hdb;
	15'h5c29: q<=8'h60;
	15'h5c2a: q<=8'had;
	15'h5c2b: q<=8'hd8;
	15'h5c2c: q<=8'h60;
	15'h5c2d: q<=8'h29;
	15'h5c2e: q<=8'h78;
	15'h5c2f: q<=8'h85;
	15'h5c30: q<=8'h4d;
	15'h5c31: q<=8'hf0;
	15'h5c32: q<=8'h05;
	15'h5c33: q<=8'h8d;
	15'h5c34: q<=8'hc0;
	15'h5c35: q<=8'h60;
	15'h5c36: q<=8'ha2;
	15'h5c37: q<=8'ha4;
	15'h5c38: q<=8'h8e;
	15'h5c39: q<=8'hc1;
	15'h5c3a: q<=8'h60;
	15'h5c3b: q<=8'ha2;
	15'h5c3c: q<=8'h00;
	15'h5c3d: q<=8'ha5;
	15'h5c3e: q<=8'h4e;
	15'h5c3f: q<=8'hf0;
	15'h5c40: q<=8'h06;
	15'h5c41: q<=8'h0a;
	15'h5c42: q<=8'h8d;
	15'h5c43: q<=8'hc2;
	15'h5c44: q<=8'h60;
	15'h5c45: q<=8'ha2;
	15'h5c46: q<=8'ha4;
	15'h5c47: q<=8'h8e;
	15'h5c48: q<=8'hc3;
	15'h5c49: q<=8'h60;
	15'h5c4a: q<=8'h20;
	15'h5c4b: q<=8'h0d;
	15'h5c4c: q<=8'hdd;
	15'h5c4d: q<=8'ha4;
	15'h5c4e: q<=8'h4d;
	15'h5c4f: q<=8'ha9;
	15'h5c50: q<=8'hd0;
	15'h5c51: q<=8'ha2;
	15'h5c52: q<=8'hf0;
	15'h5c53: q<=8'h20;
	15'h5c54: q<=8'h2b;
	15'h5c55: q<=8'hdd;
	15'h5c56: q<=8'ha4;
	15'h5c57: q<=8'h4e;
	15'h5c58: q<=8'h20;
	15'h5c59: q<=8'h27;
	15'h5c5a: q<=8'hdd;
	15'h5c5b: q<=8'ha5;
	15'h5c5c: q<=8'h52;
	15'h5c5d: q<=8'h29;
	15'h5c5e: q<=8'h10;
	15'h5c5f: q<=8'hf0;
	15'h5c60: q<=8'h1d;
	15'h5c61: q<=8'ha9;
	15'h5c62: q<=8'h34;
	15'h5c63: q<=8'ha2;
	15'h5c64: q<=8'h82;
	15'h5c65: q<=8'h20;
	15'h5c66: q<=8'h39;
	15'h5c67: q<=8'hdf;
	15'h5c68: q<=8'ha0;
	15'h5c69: q<=8'h10;
	15'h5c6a: q<=8'ha5;
	15'h5c6b: q<=8'h4d;
	15'h5c6c: q<=8'h29;
	15'h5c6d: q<=8'h60;
	15'h5c6e: q<=8'hf0;
	15'h5c6f: q<=8'h0e;
	15'h5c70: q<=8'h49;
	15'h5c71: q<=8'h20;
	15'h5c72: q<=8'hf0;
	15'h5c73: q<=8'h04;
	15'h5c74: q<=8'ha9;
	15'h5c75: q<=8'h04;
	15'h5c76: q<=8'ha0;
	15'h5c77: q<=8'h08;
	15'h5c78: q<=8'h8d;
	15'h5c79: q<=8'he0;
	15'h5c7a: q<=8'h60;
	15'h5c7b: q<=8'h8c;
	15'h5c7c: q<=8'h00;
	15'h5c7d: q<=8'h40;
	15'h5c7e: q<=8'ha9;
	15'h5c7f: q<=8'h34;
	15'h5c80: q<=8'ha2;
	15'h5c81: q<=8'h92;
	15'h5c82: q<=8'h20;
	15'h5c83: q<=8'h39;
	15'h5c84: q<=8'hdf;
	15'h5c85: q<=8'ha2;
	15'h5c86: q<=8'h0b;
	15'h5c87: q<=8'hb5;
	15'h5c88: q<=8'h7d;
	15'h5c89: q<=8'hf0;
	15'h5c8a: q<=8'h19;
	15'h5c8b: q<=8'h85;
	15'h5c8c: q<=8'h35;
	15'h5c8d: q<=8'h86;
	15'h5c8e: q<=8'h38;
	15'h5c8f: q<=8'h8a;
	15'h5c90: q<=8'h20;
	15'h5c91: q<=8'h1f;
	15'h5c92: q<=8'hdf;
	15'h5c93: q<=8'ha0;
	15'h5c94: q<=8'hf4;
	15'h5c95: q<=8'ha2;
	15'h5c96: q<=8'hf4;
	15'h5c97: q<=8'ha5;
	15'h5c98: q<=8'h35;
	15'h5c99: q<=8'h20;
	15'h5c9a: q<=8'ha9;
	15'h5c9b: q<=8'hd8;
	15'h5c9c: q<=8'ha9;
	15'h5c9d: q<=8'h0c;
	15'h5c9e: q<=8'haa;
	15'h5c9f: q<=8'h20;
	15'h5ca0: q<=8'h75;
	15'h5ca1: q<=8'hdf;
	15'h5ca2: q<=8'ha6;
	15'h5ca3: q<=8'h38;
	15'h5ca4: q<=8'hca;
	15'h5ca5: q<=8'h10;
	15'h5ca6: q<=8'he0;
	15'h5ca7: q<=8'h20;
	15'h5ca8: q<=8'h53;
	15'h5ca9: q<=8'hdf;
	15'h5caa: q<=8'ha9;
	15'h5cab: q<=8'h00;
	15'h5cac: q<=8'ha2;
	15'h5cad: q<=8'h16;
	15'h5cae: q<=8'h20;
	15'h5caf: q<=8'h75;
	15'h5cb0: q<=8'hdf;
	15'h5cb1: q<=8'ha2;
	15'h5cb2: q<=8'h04;
	15'h5cb3: q<=8'h86;
	15'h5cb4: q<=8'h37;
	15'h5cb5: q<=8'ha6;
	15'h5cb6: q<=8'h37;
	15'h5cb7: q<=8'ha0;
	15'h5cb8: q<=8'h00;
	15'h5cb9: q<=8'hb5;
	15'h5cba: q<=8'h78;
	15'h5cbb: q<=8'hf0;
	15'h5cbc: q<=8'h03;
	15'h5cbd: q<=8'hbc;
	15'h5cbe: q<=8'he1;
	15'h5cbf: q<=8'hdc;
	15'h5cc0: q<=8'hb9;
	15'h5cc1: q<=8'he4;
	15'h5cc2: q<=8'h31;
	15'h5cc3: q<=8'hbe;
	15'h5cc4: q<=8'he5;
	15'h5cc5: q<=8'h31;
	15'h5cc6: q<=8'h20;
	15'h5cc7: q<=8'h57;
	15'h5cc8: q<=8'hdf;
	15'h5cc9: q<=8'hc6;
	15'h5cca: q<=8'h37;
	15'h5ccb: q<=8'h10;
	15'h5ccc: q<=8'he8;
	15'h5ccd: q<=8'ha2;
	15'h5cce: q<=8'hac;
	15'h5ccf: q<=8'ha9;
	15'h5cd0: q<=8'h30;
	15'h5cd1: q<=8'h20;
	15'h5cd2: q<=8'h75;
	15'h5cd3: q<=8'hdf;
	15'h5cd4: q<=8'ha4;
	15'h5cd5: q<=8'h50;
	15'h5cd6: q<=8'hb9;
	15'h5cd7: q<=8'he8;
	15'h5cd8: q<=8'hdf;
	15'h5cd9: q<=8'hbe;
	15'h5cda: q<=8'he4;
	15'h5cdb: q<=8'hdf;
	15'h5cdc: q<=8'ha0;
	15'h5cdd: q<=8'hc0;
	15'h5cde: q<=8'h4c;
	15'h5cdf: q<=8'h73;
	15'h5ce0: q<=8'hdf;
	15'h5ce1: q<=8'h2e;
	15'h5ce2: q<=8'h38;
	15'h5ce3: q<=8'h34;
	15'h5ce4: q<=8'h36;
	15'h5ce5: q<=8'h1e;
	15'h5ce6: q<=8'ha0;
	15'h5ce7: q<=8'h00;
	15'h5ce8: q<=8'h84;
	15'h5ce9: q<=8'h73;
	15'h5cea: q<=8'h8c;
	15'h5ceb: q<=8'h14;
	15'h5cec: q<=8'h04;
	15'h5ced: q<=8'h8d;
	15'h5cee: q<=8'h8e;
	15'h5cef: q<=8'h60;
	15'h5cf0: q<=8'h8e;
	15'h5cf1: q<=8'h8f;
	15'h5cf2: q<=8'h60;
	15'h5cf3: q<=8'h8c;
	15'h5cf4: q<=8'h90;
	15'h5cf5: q<=8'h60;
	15'h5cf6: q<=8'ha2;
	15'h5cf7: q<=8'h10;
	15'h5cf8: q<=8'h8e;
	15'h5cf9: q<=8'h8c;
	15'h5cfa: q<=8'h60;
	15'h5cfb: q<=8'h8e;
	15'h5cfc: q<=8'h94;
	15'h5cfd: q<=8'h60;
	15'h5cfe: q<=8'hca;
	15'h5cff: q<=8'h30;
	15'h5d00: q<=8'h0b;
	15'h5d01: q<=8'had;
	15'h5d02: q<=8'h40;
	15'h5d03: q<=8'h60;
	15'h5d04: q<=8'h30;
	15'h5d05: q<=8'hf8;
	15'h5d06: q<=8'had;
	15'h5d07: q<=8'h60;
	15'h5d08: q<=8'h60;
	15'h5d09: q<=8'hac;
	15'h5d0a: q<=8'h70;
	15'h5d0b: q<=8'h60;
	15'h5d0c: q<=8'h60;
	15'h5d0d: q<=8'h20;
	15'h5d0e: q<=8'h53;
	15'h5d0f: q<=8'hdf;
	15'h5d10: q<=8'ha9;
	15'h5d11: q<=8'h00;
	15'h5d12: q<=8'h20;
	15'h5d13: q<=8'h6a;
	15'h5d14: q<=8'hdf;
	15'h5d15: q<=8'ha9;
	15'h5d16: q<=8'he8;
	15'h5d17: q<=8'hac;
	15'h5d18: q<=8'h00;
	15'h5d19: q<=8'h0d;
	15'h5d1a: q<=8'h20;
	15'h5d1b: q<=8'h29;
	15'h5d1c: q<=8'hdd;
	15'h5d1d: q<=8'hac;
	15'h5d1e: q<=8'h00;
	15'h5d1f: q<=8'h0e;
	15'h5d20: q<=8'h20;
	15'h5d21: q<=8'h27;
	15'h5d22: q<=8'hdd;
	15'h5d23: q<=8'h20;
	15'h5d24: q<=8'he0;
	15'h5d25: q<=8'hdb;
	15'h5d26: q<=8'ha8;
	15'h5d27: q<=8'ha9;
	15'h5d28: q<=8'hd0;
	15'h5d29: q<=8'ha2;
	15'h5d2a: q<=8'hf8;
	15'h5d2b: q<=8'h84;
	15'h5d2c: q<=8'h35;
	15'h5d2d: q<=8'h20;
	15'h5d2e: q<=8'h75;
	15'h5d2f: q<=8'hdf;
	15'h5d30: q<=8'ha2;
	15'h5d31: q<=8'h07;
	15'h5d32: q<=8'h86;
	15'h5d33: q<=8'h37;
	15'h5d34: q<=8'h06;
	15'h5d35: q<=8'h35;
	15'h5d36: q<=8'ha9;
	15'h5d37: q<=8'h00;
	15'h5d38: q<=8'h2a;
	15'h5d39: q<=8'h20;
	15'h5d3a: q<=8'h1f;
	15'h5d3b: q<=8'hdf;
	15'h5d3c: q<=8'hc6;
	15'h5d3d: q<=8'h37;
	15'h5d3e: q<=8'h10;
	15'h5d3f: q<=8'hf4;
	15'h5d40: q<=8'h60;
	15'h5d41: q<=8'had;
	15'h5d42: q<=8'h0f;
	15'h5d43: q<=8'h04;
	15'h5d44: q<=8'h0a;
	15'h5d45: q<=8'h85;
	15'h5d46: q<=8'h29;
	15'h5d47: q<=8'had;
	15'h5d48: q<=8'h10;
	15'h5d49: q<=8'h04;
	15'h5d4a: q<=8'h2a;
	15'h5d4b: q<=8'h85;
	15'h5d4c: q<=8'h2a;
	15'h5d4d: q<=8'had;
	15'h5d4e: q<=8'h0c;
	15'h5d4f: q<=8'h04;
	15'h5d50: q<=8'h18;
	15'h5d51: q<=8'h65;
	15'h5d52: q<=8'h29;
	15'h5d53: q<=8'h8d;
	15'h5d54: q<=8'h95;
	15'h5d55: q<=8'h60;
	15'h5d56: q<=8'h85;
	15'h5d57: q<=8'h29;
	15'h5d58: q<=8'had;
	15'h5d59: q<=8'h0d;
	15'h5d5a: q<=8'h04;
	15'h5d5b: q<=8'h65;
	15'h5d5c: q<=8'h2a;
	15'h5d5d: q<=8'h8d;
	15'h5d5e: q<=8'h96;
	15'h5d5f: q<=8'h60;
	15'h5d60: q<=8'h05;
	15'h5d61: q<=8'h29;
	15'h5d62: q<=8'hd0;
	15'h5d63: q<=8'h05;
	15'h5d64: q<=8'ha9;
	15'h5d65: q<=8'h01;
	15'h5d66: q<=8'h8d;
	15'h5d67: q<=8'h95;
	15'h5d68: q<=8'h60;
	15'h5d69: q<=8'had;
	15'h5d6a: q<=8'h09;
	15'h5d6b: q<=8'h04;
	15'h5d6c: q<=8'h8d;
	15'h5d6d: q<=8'h8d;
	15'h5d6e: q<=8'h60;
	15'h5d6f: q<=8'had;
	15'h5d70: q<=8'h0a;
	15'h5d71: q<=8'h04;
	15'h5d72: q<=8'hae;
	15'h5d73: q<=8'h0b;
	15'h5d74: q<=8'h04;
	15'h5d75: q<=8'h20;
	15'h5d76: q<=8'he6;
	15'h5d77: q<=8'hdc;
	15'h5d78: q<=8'h8d;
	15'h5d79: q<=8'h12;
	15'h5d7a: q<=8'h04;
	15'h5d7b: q<=8'h8c;
	15'h5d7c: q<=8'h13;
	15'h5d7d: q<=8'h04;
	15'h5d7e: q<=8'ha9;
	15'h5d7f: q<=8'h3d;
	15'h5d80: q<=8'ha2;
	15'h5d81: q<=8'hce;
	15'h5d82: q<=8'h20;
	15'h5d83: q<=8'h39;
	15'h5d84: q<=8'hdf;
	15'h5d85: q<=8'ha9;
	15'h5d86: q<=8'h06;
	15'h5d87: q<=8'h85;
	15'h5d88: q<=8'h3b;
	15'h5d89: q<=8'ha9;
	15'h5d8a: q<=8'h04;
	15'h5d8b: q<=8'h85;
	15'h5d8c: q<=8'h3c;
	15'h5d8d: q<=8'h85;
	15'h5d8e: q<=8'h37;
	15'h5d8f: q<=8'ha0;
	15'h5d90: q<=8'h00;
	15'h5d91: q<=8'h84;
	15'h5d92: q<=8'h31;
	15'h5d93: q<=8'h84;
	15'h5d94: q<=8'h32;
	15'h5d95: q<=8'h84;
	15'h5d96: q<=8'h33;
	15'h5d97: q<=8'h84;
	15'h5d98: q<=8'h34;
	15'h5d99: q<=8'hb1;
	15'h5d9a: q<=8'h3b;
	15'h5d9b: q<=8'h85;
	15'h5d9c: q<=8'h56;
	15'h5d9d: q<=8'he6;
	15'h5d9e: q<=8'h3b;
	15'h5d9f: q<=8'hb1;
	15'h5da0: q<=8'h3b;
	15'h5da1: q<=8'h85;
	15'h5da2: q<=8'h57;
	15'h5da3: q<=8'he6;
	15'h5da4: q<=8'h3b;
	15'h5da5: q<=8'hb1;
	15'h5da6: q<=8'h3b;
	15'h5da7: q<=8'h85;
	15'h5da8: q<=8'h58;
	15'h5da9: q<=8'he6;
	15'h5daa: q<=8'h3b;
	15'h5dab: q<=8'hf8;
	15'h5dac: q<=8'ha0;
	15'h5dad: q<=8'h17;
	15'h5dae: q<=8'h84;
	15'h5daf: q<=8'h38;
	15'h5db0: q<=8'h26;
	15'h5db1: q<=8'h56;
	15'h5db2: q<=8'h26;
	15'h5db3: q<=8'h57;
	15'h5db4: q<=8'h26;
	15'h5db5: q<=8'h58;
	15'h5db6: q<=8'ha0;
	15'h5db7: q<=8'h03;
	15'h5db8: q<=8'ha2;
	15'h5db9: q<=8'h00;
	15'h5dba: q<=8'hb5;
	15'h5dbb: q<=8'h31;
	15'h5dbc: q<=8'h75;
	15'h5dbd: q<=8'h31;
	15'h5dbe: q<=8'h95;
	15'h5dbf: q<=8'h31;
	15'h5dc0: q<=8'he8;
	15'h5dc1: q<=8'h88;
	15'h5dc2: q<=8'h10;
	15'h5dc3: q<=8'hf6;
	15'h5dc4: q<=8'hc6;
	15'h5dc5: q<=8'h38;
	15'h5dc6: q<=8'h10;
	15'h5dc7: q<=8'he8;
	15'h5dc8: q<=8'hd8;
	15'h5dc9: q<=8'ha9;
	15'h5dca: q<=8'h31;
	15'h5dcb: q<=8'ha0;
	15'h5dcc: q<=8'h04;
	15'h5dcd: q<=8'h20;
	15'h5dce: q<=8'hb1;
	15'h5dcf: q<=8'hdf;
	15'h5dd0: q<=8'ha9;
	15'h5dd1: q<=8'hd0;
	15'h5dd2: q<=8'ha2;
	15'h5dd3: q<=8'hf8;
	15'h5dd4: q<=8'h20;
	15'h5dd5: q<=8'h75;
	15'h5dd6: q<=8'hdf;
	15'h5dd7: q<=8'hc6;
	15'h5dd8: q<=8'h37;
	15'h5dd9: q<=8'h10;
	15'h5dda: q<=8'hb4;
	15'h5ddb: q<=8'h60;
	15'h5ddc: q<=8'h73;
	15'h5ddd: q<=8'h00;
	15'h5dde: q<=8'h09;
	15'h5ddf: q<=8'h0a;
	15'h5de0: q<=8'h15;
	15'h5de1: q<=8'h16;
	15'h5de2: q<=8'h22;
	15'h5de3: q<=8'h15;
	15'h5de4: q<=8'h06;
	15'h5de5: q<=8'h15;
	15'h5de6: q<=8'h07;
	15'h5de7: q<=8'h06;
	15'h5de8: q<=8'h04;
	15'h5de9: q<=8'ha9;
	15'h5dea: q<=8'h04;
	15'h5deb: q<=8'hd0;
	15'h5dec: q<=8'h06;
	15'h5ded: q<=8'ha9;
	15'h5dee: q<=8'h03;
	15'h5def: q<=8'hd0;
	15'h5df0: q<=8'h02;
	15'h5df1: q<=8'ha9;
	15'h5df2: q<=8'h07;
	15'h5df3: q<=8'ha0;
	15'h5df4: q<=8'hff;
	15'h5df5: q<=8'hd0;
	15'h5df6: q<=8'h08;
	15'h5df7: q<=8'ha9;
	15'h5df8: q<=8'h03;
	15'h5df9: q<=8'hd0;
	15'h5dfa: q<=8'h02;
	15'h5dfb: q<=8'ha9;
	15'h5dfc: q<=8'h04;
	15'h5dfd: q<=8'ha0;
	15'h5dfe: q<=8'h00;
	15'h5dff: q<=8'h8c;
	15'h5e00: q<=8'hc6;
	15'h5e01: q<=8'h01;
	15'h5e02: q<=8'h48;
	15'h5e03: q<=8'h0d;
	15'h5e04: q<=8'hc7;
	15'h5e05: q<=8'h01;
	15'h5e06: q<=8'h8d;
	15'h5e07: q<=8'hc7;
	15'h5e08: q<=8'h01;
	15'h5e09: q<=8'h68;
	15'h5e0a: q<=8'h0d;
	15'h5e0b: q<=8'hc8;
	15'h5e0c: q<=8'h01;
	15'h5e0d: q<=8'h8d;
	15'h5e0e: q<=8'hc8;
	15'h5e0f: q<=8'h01;
	15'h5e10: q<=8'h60;
	15'h5e11: q<=8'ha9;
	15'h5e12: q<=8'h07;
	15'h5e13: q<=8'h8d;
	15'h5e14: q<=8'hc7;
	15'h5e15: q<=8'h01;
	15'h5e16: q<=8'ha9;
	15'h5e17: q<=8'h00;
	15'h5e18: q<=8'h8d;
	15'h5e19: q<=8'hc8;
	15'h5e1a: q<=8'h01;
	15'h5e1b: q<=8'had;
	15'h5e1c: q<=8'hca;
	15'h5e1d: q<=8'h01;
	15'h5e1e: q<=8'hd0;
	15'h5e1f: q<=8'h4b;
	15'h5e20: q<=8'had;
	15'h5e21: q<=8'hc7;
	15'h5e22: q<=8'h01;
	15'h5e23: q<=8'hf0;
	15'h5e24: q<=8'h46;
	15'h5e25: q<=8'ha2;
	15'h5e26: q<=8'h00;
	15'h5e27: q<=8'h8e;
	15'h5e28: q<=8'hcb;
	15'h5e29: q<=8'h01;
	15'h5e2a: q<=8'h8e;
	15'h5e2b: q<=8'hcf;
	15'h5e2c: q<=8'h01;
	15'h5e2d: q<=8'h8e;
	15'h5e2e: q<=8'hce;
	15'h5e2f: q<=8'h01;
	15'h5e30: q<=8'ha2;
	15'h5e31: q<=8'h08;
	15'h5e32: q<=8'h38;
	15'h5e33: q<=8'h6e;
	15'h5e34: q<=8'hce;
	15'h5e35: q<=8'h01;
	15'h5e36: q<=8'h0a;
	15'h5e37: q<=8'hca;
	15'h5e38: q<=8'h90;
	15'h5e39: q<=8'hf9;
	15'h5e3a: q<=8'ha0;
	15'h5e3b: q<=8'h80;
	15'h5e3c: q<=8'had;
	15'h5e3d: q<=8'hce;
	15'h5e3e: q<=8'h01;
	15'h5e3f: q<=8'h2d;
	15'h5e40: q<=8'hc8;
	15'h5e41: q<=8'h01;
	15'h5e42: q<=8'hd0;
	15'h5e43: q<=8'h02;
	15'h5e44: q<=8'ha0;
	15'h5e45: q<=8'h20;
	15'h5e46: q<=8'h8c;
	15'h5e47: q<=8'hca;
	15'h5e48: q<=8'h01;
	15'h5e49: q<=8'had;
	15'h5e4a: q<=8'hce;
	15'h5e4b: q<=8'h01;
	15'h5e4c: q<=8'h4d;
	15'h5e4d: q<=8'hc7;
	15'h5e4e: q<=8'h01;
	15'h5e4f: q<=8'h8d;
	15'h5e50: q<=8'hc7;
	15'h5e51: q<=8'h01;
	15'h5e52: q<=8'h8a;
	15'h5e53: q<=8'h0a;
	15'h5e54: q<=8'haa;
	15'h5e55: q<=8'hbd;
	15'h5e56: q<=8'hdd;
	15'h5e57: q<=8'hdd;
	15'h5e58: q<=8'h8d;
	15'h5e59: q<=8'hcc;
	15'h5e5a: q<=8'h01;
	15'h5e5b: q<=8'hbd;
	15'h5e5c: q<=8'hde;
	15'h5e5d: q<=8'hdd;
	15'h5e5e: q<=8'h8d;
	15'h5e5f: q<=8'hcd;
	15'h5e60: q<=8'h01;
	15'h5e61: q<=8'hbd;
	15'h5e62: q<=8'he3;
	15'h5e63: q<=8'hdd;
	15'h5e64: q<=8'h85;
	15'h5e65: q<=8'hbd;
	15'h5e66: q<=8'hbd;
	15'h5e67: q<=8'he4;
	15'h5e68: q<=8'hdd;
	15'h5e69: q<=8'h85;
	15'h5e6a: q<=8'hbe;
	15'h5e6b: q<=8'ha0;
	15'h5e6c: q<=8'h00;
	15'h5e6d: q<=8'h8c;
	15'h5e6e: q<=8'h40;
	15'h5e6f: q<=8'h60;
	15'h5e70: q<=8'had;
	15'h5e71: q<=8'hca;
	15'h5e72: q<=8'h01;
	15'h5e73: q<=8'hd0;
	15'h5e74: q<=8'h01;
	15'h5e75: q<=8'h60;
	15'h5e76: q<=8'hac;
	15'h5e77: q<=8'hcb;
	15'h5e78: q<=8'h01;
	15'h5e79: q<=8'hae;
	15'h5e7a: q<=8'hcc;
	15'h5e7b: q<=8'h01;
	15'h5e7c: q<=8'h0a;
	15'h5e7d: q<=8'h90;
	15'h5e7e: q<=8'h0d;
	15'h5e7f: q<=8'h9d;
	15'h5e80: q<=8'h00;
	15'h5e81: q<=8'h60;
	15'h5e82: q<=8'ha9;
	15'h5e83: q<=8'h40;
	15'h5e84: q<=8'h8d;
	15'h5e85: q<=8'hca;
	15'h5e86: q<=8'h01;
	15'h5e87: q<=8'ha0;
	15'h5e88: q<=8'h0e;
	15'h5e89: q<=8'hb8;
	15'h5e8a: q<=8'h50;
	15'h5e8b: q<=8'h73;
	15'h5e8c: q<=8'h10;
	15'h5e8d: q<=8'h25;
	15'h5e8e: q<=8'ha9;
	15'h5e8f: q<=8'h80;
	15'h5e90: q<=8'h8d;
	15'h5e91: q<=8'hca;
	15'h5e92: q<=8'h01;
	15'h5e93: q<=8'had;
	15'h5e94: q<=8'hc6;
	15'h5e95: q<=8'h01;
	15'h5e96: q<=8'hf0;
	15'h5e97: q<=8'h04;
	15'h5e98: q<=8'ha9;
	15'h5e99: q<=8'h00;
	15'h5e9a: q<=8'h91;
	15'h5e9b: q<=8'hbd;
	15'h5e9c: q<=8'hb1;
	15'h5e9d: q<=8'hbd;
	15'h5e9e: q<=8'hec;
	15'h5e9f: q<=8'hcd;
	15'h5ea0: q<=8'h01;
	15'h5ea1: q<=8'h90;
	15'h5ea2: q<=8'h08;
	15'h5ea3: q<=8'ha9;
	15'h5ea4: q<=8'h00;
	15'h5ea5: q<=8'h8d;
	15'h5ea6: q<=8'hca;
	15'h5ea7: q<=8'h01;
	15'h5ea8: q<=8'had;
	15'h5ea9: q<=8'hcf;
	15'h5eaa: q<=8'h01;
	15'h5eab: q<=8'h9d;
	15'h5eac: q<=8'h00;
	15'h5ead: q<=8'h60;
	15'h5eae: q<=8'ha0;
	15'h5eaf: q<=8'h0c;
	15'h5eb0: q<=8'hb8;
	15'h5eb1: q<=8'h50;
	15'h5eb2: q<=8'h3f;
	15'h5eb3: q<=8'ha9;
	15'h5eb4: q<=8'h08;
	15'h5eb5: q<=8'h8d;
	15'h5eb6: q<=8'h40;
	15'h5eb7: q<=8'h60;
	15'h5eb8: q<=8'h9d;
	15'h5eb9: q<=8'h00;
	15'h5eba: q<=8'h60;
	15'h5ebb: q<=8'ha9;
	15'h5ebc: q<=8'h09;
	15'h5ebd: q<=8'h8d;
	15'h5ebe: q<=8'h40;
	15'h5ebf: q<=8'h60;
	15'h5ec0: q<=8'hea;
	15'h5ec1: q<=8'ha9;
	15'h5ec2: q<=8'h08;
	15'h5ec3: q<=8'h8d;
	15'h5ec4: q<=8'h40;
	15'h5ec5: q<=8'h60;
	15'h5ec6: q<=8'hec;
	15'h5ec7: q<=8'hcd;
	15'h5ec8: q<=8'h01;
	15'h5ec9: q<=8'had;
	15'h5eca: q<=8'h50;
	15'h5ecb: q<=8'h60;
	15'h5ecc: q<=8'h90;
	15'h5ecd: q<=8'h20;
	15'h5ece: q<=8'h4d;
	15'h5ecf: q<=8'hcf;
	15'h5ed0: q<=8'h01;
	15'h5ed1: q<=8'hf0;
	15'h5ed2: q<=8'h13;
	15'h5ed3: q<=8'ha9;
	15'h5ed4: q<=8'h00;
	15'h5ed5: q<=8'hac;
	15'h5ed6: q<=8'hcb;
	15'h5ed7: q<=8'h01;
	15'h5ed8: q<=8'h91;
	15'h5ed9: q<=8'hbd;
	15'h5eda: q<=8'h88;
	15'h5edb: q<=8'h10;
	15'h5edc: q<=8'hfb;
	15'h5edd: q<=8'had;
	15'h5ede: q<=8'hce;
	15'h5edf: q<=8'h01;
	15'h5ee0: q<=8'h0d;
	15'h5ee1: q<=8'hc9;
	15'h5ee2: q<=8'h01;
	15'h5ee3: q<=8'h8d;
	15'h5ee4: q<=8'hc9;
	15'h5ee5: q<=8'h01;
	15'h5ee6: q<=8'ha9;
	15'h5ee7: q<=8'h00;
	15'h5ee8: q<=8'h8d;
	15'h5ee9: q<=8'hca;
	15'h5eea: q<=8'h01;
	15'h5eeb: q<=8'hb8;
	15'h5eec: q<=8'h50;
	15'h5eed: q<=8'h02;
	15'h5eee: q<=8'h91;
	15'h5eef: q<=8'hbd;
	15'h5ef0: q<=8'ha0;
	15'h5ef1: q<=8'h00;
	15'h5ef2: q<=8'h18;
	15'h5ef3: q<=8'h6d;
	15'h5ef4: q<=8'hcf;
	15'h5ef5: q<=8'h01;
	15'h5ef6: q<=8'h8d;
	15'h5ef7: q<=8'hcf;
	15'h5ef8: q<=8'h01;
	15'h5ef9: q<=8'hee;
	15'h5efa: q<=8'hcb;
	15'h5efb: q<=8'h01;
	15'h5efc: q<=8'hee;
	15'h5efd: q<=8'hcc;
	15'h5efe: q<=8'h01;
	15'h5eff: q<=8'h8c;
	15'h5f00: q<=8'h40;
	15'h5f01: q<=8'h60;
	15'h5f02: q<=8'h98;
	15'h5f03: q<=8'hd0;
	15'h5f04: q<=8'h03;
	15'h5f05: q<=8'h4c;
	15'h5f06: q<=8'h1b;
	15'h5f07: q<=8'hde;
	15'h5f08: q<=8'h60;
	15'h5f09: q<=8'ha9;
	15'h5f0a: q<=8'hc0;
	15'h5f0b: q<=8'hd0;
	15'h5f0c: q<=8'h05;
	15'h5f0d: q<=8'h20;
	15'h5f0e: q<=8'h53;
	15'h5f0f: q<=8'hdf;
	15'h5f10: q<=8'ha9;
	15'h5f11: q<=8'h20;
	15'h5f12: q<=8'ha0;
	15'h5f13: q<=8'h00;
	15'h5f14: q<=8'h91;
	15'h5f15: q<=8'h74;
	15'h5f16: q<=8'h4c;
	15'h5f17: q<=8'hac;
	15'h5f18: q<=8'hdf;
	15'h5f19: q<=8'h90;
	15'h5f1a: q<=8'h04;
	15'h5f1b: q<=8'h29;
	15'h5f1c: q<=8'h0f;
	15'h5f1d: q<=8'hf0;
	15'h5f1e: q<=8'h05;
	15'h5f1f: q<=8'h29;
	15'h5f20: q<=8'h0f;
	15'h5f21: q<=8'h18;
	15'h5f22: q<=8'h69;
	15'h5f23: q<=8'h01;
	15'h5f24: q<=8'h08;
	15'h5f25: q<=8'h0a;
	15'h5f26: q<=8'ha0;
	15'h5f27: q<=8'h00;
	15'h5f28: q<=8'haa;
	15'h5f29: q<=8'hbd;
	15'h5f2a: q<=8'he4;
	15'h5f2b: q<=8'h31;
	15'h5f2c: q<=8'h91;
	15'h5f2d: q<=8'h74;
	15'h5f2e: q<=8'hbd;
	15'h5f2f: q<=8'he5;
	15'h5f30: q<=8'h31;
	15'h5f31: q<=8'hc8;
	15'h5f32: q<=8'h91;
	15'h5f33: q<=8'h74;
	15'h5f34: q<=8'h20;
	15'h5f35: q<=8'h5f;
	15'h5f36: q<=8'hdf;
	15'h5f37: q<=8'h28;
	15'h5f38: q<=8'h60;
	15'h5f39: q<=8'h4a;
	15'h5f3a: q<=8'h29;
	15'h5f3b: q<=8'h0f;
	15'h5f3c: q<=8'h09;
	15'h5f3d: q<=8'ha0;
	15'h5f3e: q<=8'ha0;
	15'h5f3f: q<=8'h01;
	15'h5f40: q<=8'h91;
	15'h5f41: q<=8'h74;
	15'h5f42: q<=8'h88;
	15'h5f43: q<=8'h8a;
	15'h5f44: q<=8'h6a;
	15'h5f45: q<=8'h91;
	15'h5f46: q<=8'h74;
	15'h5f47: q<=8'hc8;
	15'h5f48: q<=8'hd0;
	15'h5f49: q<=8'h15;
	15'h5f4a: q<=8'ha4;
	15'h5f4b: q<=8'h73;
	15'h5f4c: q<=8'h09;
	15'h5f4d: q<=8'h60;
	15'h5f4e: q<=8'haa;
	15'h5f4f: q<=8'h98;
	15'h5f50: q<=8'h4c;
	15'h5f51: q<=8'h57;
	15'h5f52: q<=8'hdf;
	15'h5f53: q<=8'ha9;
	15'h5f54: q<=8'h40;
	15'h5f55: q<=8'ha2;
	15'h5f56: q<=8'h80;
	15'h5f57: q<=8'ha0;
	15'h5f58: q<=8'h00;
	15'h5f59: q<=8'h91;
	15'h5f5a: q<=8'h74;
	15'h5f5b: q<=8'hc8;
	15'h5f5c: q<=8'h8a;
	15'h5f5d: q<=8'h91;
	15'h5f5e: q<=8'h74;
	15'h5f5f: q<=8'h98;
	15'h5f60: q<=8'h38;
	15'h5f61: q<=8'h65;
	15'h5f62: q<=8'h74;
	15'h5f63: q<=8'h85;
	15'h5f64: q<=8'h74;
	15'h5f65: q<=8'h90;
	15'h5f66: q<=8'h02;
	15'h5f67: q<=8'he6;
	15'h5f68: q<=8'h75;
	15'h5f69: q<=8'h60;
	15'h5f6a: q<=8'ha0;
	15'h5f6b: q<=8'h00;
	15'h5f6c: q<=8'h09;
	15'h5f6d: q<=8'h70;
	15'h5f6e: q<=8'haa;
	15'h5f6f: q<=8'h98;
	15'h5f70: q<=8'h4c;
	15'h5f71: q<=8'h57;
	15'h5f72: q<=8'hdf;
	15'h5f73: q<=8'h84;
	15'h5f74: q<=8'h73;
	15'h5f75: q<=8'ha0;
	15'h5f76: q<=8'h00;
	15'h5f77: q<=8'h0a;
	15'h5f78: q<=8'h90;
	15'h5f79: q<=8'h01;
	15'h5f7a: q<=8'h88;
	15'h5f7b: q<=8'h84;
	15'h5f7c: q<=8'h6f;
	15'h5f7d: q<=8'h0a;
	15'h5f7e: q<=8'h26;
	15'h5f7f: q<=8'h6f;
	15'h5f80: q<=8'h85;
	15'h5f81: q<=8'h6e;
	15'h5f82: q<=8'h8a;
	15'h5f83: q<=8'h0a;
	15'h5f84: q<=8'ha0;
	15'h5f85: q<=8'h00;
	15'h5f86: q<=8'h90;
	15'h5f87: q<=8'h01;
	15'h5f88: q<=8'h88;
	15'h5f89: q<=8'h84;
	15'h5f8a: q<=8'h71;
	15'h5f8b: q<=8'h0a;
	15'h5f8c: q<=8'h26;
	15'h5f8d: q<=8'h71;
	15'h5f8e: q<=8'h85;
	15'h5f8f: q<=8'h70;
	15'h5f90: q<=8'ha2;
	15'h5f91: q<=8'h6e;
	15'h5f92: q<=8'ha0;
	15'h5f93: q<=8'h00;
	15'h5f94: q<=8'hb5;
	15'h5f95: q<=8'h02;
	15'h5f96: q<=8'h91;
	15'h5f97: q<=8'h74;
	15'h5f98: q<=8'hb5;
	15'h5f99: q<=8'h03;
	15'h5f9a: q<=8'h29;
	15'h5f9b: q<=8'h1f;
	15'h5f9c: q<=8'hc8;
	15'h5f9d: q<=8'h91;
	15'h5f9e: q<=8'h74;
	15'h5f9f: q<=8'hb5;
	15'h5fa0: q<=8'h00;
	15'h5fa1: q<=8'hc8;
	15'h5fa2: q<=8'h91;
	15'h5fa3: q<=8'h74;
	15'h5fa4: q<=8'hb5;
	15'h5fa5: q<=8'h01;
	15'h5fa6: q<=8'h45;
	15'h5fa7: q<=8'h73;
	15'h5fa8: q<=8'h29;
	15'h5fa9: q<=8'h1f;
	15'h5faa: q<=8'h45;
	15'h5fab: q<=8'h73;
	15'h5fac: q<=8'hc8;
	15'h5fad: q<=8'h91;
	15'h5fae: q<=8'h74;
	15'h5faf: q<=8'hd0;
	15'h5fb0: q<=8'hae;
	15'h5fb1: q<=8'h38;
	15'h5fb2: q<=8'h08;
	15'h5fb3: q<=8'h88;
	15'h5fb4: q<=8'h84;
	15'h5fb5: q<=8'hae;
	15'h5fb6: q<=8'h18;
	15'h5fb7: q<=8'h65;
	15'h5fb8: q<=8'hae;
	15'h5fb9: q<=8'h28;
	15'h5fba: q<=8'haa;
	15'h5fbb: q<=8'h08;
	15'h5fbc: q<=8'h86;
	15'h5fbd: q<=8'haf;
	15'h5fbe: q<=8'hb5;
	15'h5fbf: q<=8'h00;
	15'h5fc0: q<=8'h4a;
	15'h5fc1: q<=8'h4a;
	15'h5fc2: q<=8'h4a;
	15'h5fc3: q<=8'h4a;
	15'h5fc4: q<=8'h28;
	15'h5fc5: q<=8'h20;
	15'h5fc6: q<=8'h19;
	15'h5fc7: q<=8'hdf;
	15'h5fc8: q<=8'ha5;
	15'h5fc9: q<=8'hae;
	15'h5fca: q<=8'hd0;
	15'h5fcb: q<=8'h01;
	15'h5fcc: q<=8'h18;
	15'h5fcd: q<=8'ha6;
	15'h5fce: q<=8'haf;
	15'h5fcf: q<=8'hb5;
	15'h5fd0: q<=8'h00;
	15'h5fd1: q<=8'h20;
	15'h5fd2: q<=8'h19;
	15'h5fd3: q<=8'hdf;
	15'h5fd4: q<=8'ha6;
	15'h5fd5: q<=8'haf;
	15'h5fd6: q<=8'hca;
	15'h5fd7: q<=8'hc6;
	15'h5fd8: q<=8'hae;
	15'h5fd9: q<=8'h10;
	15'h5fda: q<=8'he0;
	15'h5fdb: q<=8'h60;
	15'h5fdc: q<=8'h10;
	15'h5fdd: q<=8'h10;
	15'h5fde: q<=8'h40;
	15'h5fdf: q<=8'h40;
	15'h5fe0: q<=8'h90;
	15'h5fe1: q<=8'h90;
	15'h5fe2: q<=8'hff;
	15'h5fe3: q<=8'hff;
	15'h5fe4: q<=8'h00;
	15'h5fe5: q<=8'h0c;
	15'h5fe6: q<=8'h16;
	15'h5fe7: q<=8'h1e;
	15'h5fe8: q<=8'h20;
	15'h5fe9: q<=8'h1e;
	15'h5fea: q<=8'h16;
	15'h5feb: q<=8'h0c;
	15'h5fec: q<=8'h00;
	15'h5fed: q<=8'hf4;
	15'h5fee: q<=8'hea;
	15'h5fef: q<=8'he2;
	15'h5ff0: q<=8'he0;
	15'h5ff1: q<=8'he2;
	15'h5ff2: q<=8'hea;
	15'h5ff3: q<=8'hf4;
	15'h5ff4: q<=8'h00;
	15'h5ff5: q<=8'h0c;
	15'h5ff6: q<=8'h16;
	15'h5ff7: q<=8'h1e;
	15'h5ff8: q<=8'h00;
	15'h5ff9: q<=8'h00;
	15'h5ffa: q<=8'h04;
	15'h5ffb: q<=8'hd7;
	15'h5ffc: q<=8'h3f;
	15'h5ffd: q<=8'hd9;
	15'h5ffe: q<=8'h04;
	15'h5fff: q<=8'hd7;
	15'h6000: q<=8'he6;
	15'h6001: q<=8'h06;
	15'h6002: q<=8'h85;
	15'h6003: q<=8'h17;
	15'h6004: q<=8'ha5;
	15'h6005: q<=8'h07;
	15'h6006: q<=8'h4a;
	15'h6007: q<=8'hb0;
	15'h6008: q<=8'h27;
	15'h6009: q<=8'ha0;
	15'h600a: q<=8'h00;
	15'h600b: q<=8'ha2;
	15'h600c: q<=8'h02;
	15'h600d: q<=8'hb5;
	15'h600e: q<=8'h13;
	15'h600f: q<=8'hf0;
	15'h6010: q<=8'h09;
	15'h6011: q<=8'hc9;
	15'h6012: q<=8'h10;
	15'h6013: q<=8'h90;
	15'h6014: q<=8'h05;
	15'h6015: q<=8'h69;
	15'h6016: q<=8'hef;
	15'h6017: q<=8'hc8;
	15'h6018: q<=8'h95;
	15'h6019: q<=8'h13;
	15'h601a: q<=8'hca;
	15'h601b: q<=8'h10;
	15'h601c: q<=8'hf0;
	15'h601d: q<=8'h98;
	15'h601e: q<=8'hd0;
	15'h601f: q<=8'h10;
	15'h6020: q<=8'ha2;
	15'h6021: q<=8'h02;
	15'h6022: q<=8'hb5;
	15'h6023: q<=8'h13;
	15'h6024: q<=8'hf0;
	15'h6025: q<=8'h07;
	15'h6026: q<=8'h18;
	15'h6027: q<=8'h69;
	15'h6028: q<=8'hef;
	15'h6029: q<=8'h95;
	15'h602a: q<=8'h13;
	15'h602b: q<=8'h30;
	15'h602c: q<=8'h03;
	15'h602d: q<=8'hca;
	15'h602e: q<=8'h10;
	15'h602f: q<=8'hf2;
	15'h6030: q<=8'h60;
	15'h6031: q<=8'h5d;
	15'h6032: q<=8'hd1;
	15'h6033: q<=8'h8f;
	15'h6034: q<=8'hd1;
	15'h6035: q<=8'h8f;
	15'h6036: q<=8'hd1;
	15'h6037: q<=8'hb1;
	15'h6038: q<=8'hd1;
	15'h6039: q<=8'heb;
	15'h603a: q<=8'hd1;
	15'h603b: q<=8'h03;
	15'h603c: q<=8'hd2;
	15'h603d: q<=8'h61;
	15'h603e: q<=8'hd2;
	15'h603f: q<=8'hcb;
	15'h6040: q<=8'hd2;
	15'h6041: q<=8'h33;
	15'h6042: q<=8'hd3;
	15'h6043: q<=8'h66;
	15'h6044: q<=8'hd3;
	15'h6045: q<=8'hb0;
	15'h6046: q<=8'hd3;
	15'h6047: q<=8'he6;
	15'h6048: q<=8'hd3;
	15'h6049: q<=8'hff;
	15'h604a: q<=8'hd3;
	15'h604b: q<=8'h17;
	15'h604c: q<=8'hd4;
	15'h604d: q<=8'h1d;
	15'h604e: q<=8'hd4;
	15'h604f: q<=8'h34;
	15'h6050: q<=8'hd4;
	15'h6051: q<=8'h4c;
	15'h6052: q<=8'hd4;
	15'h6053: q<=8'h60;
	15'h6054: q<=8'hd4;
	15'h6055: q<=8'ha1;
	15'h6056: q<=8'hd4;
	15'h6057: q<=8'hab;
	15'h6058: q<=8'hd4;
	15'h6059: q<=8'hef;
	15'h605a: q<=8'hd4;
	15'h605b: q<=8'h30;
	15'h605c: q<=8'hd5;
	15'h605d: q<=8'h75;
	15'h605e: q<=8'hd5;
	15'h605f: q<=8'h85;
	15'h6060: q<=8'hd5;
	15'h6061: q<=8'ha1;
	15'h6062: q<=8'hd5;
	15'h6063: q<=8'ha8;
	15'h6064: q<=8'hd5;
	15'h6065: q<=8'he9;
	15'h6066: q<=8'hd5;
	15'h6067: q<=8'h1c;
	15'h6068: q<=8'hd6;
	15'h6069: q<=8'h62;
	15'h606a: q<=8'hd6;
	15'h606b: q<=8'h7a;
	15'h606c: q<=8'hd6;
	15'h606d: q<=8'h67;
	15'h606e: q<=8'hd1;
	15'h606f: q<=8'h97;
	15'h6070: q<=8'hd1;
	15'h6071: q<=8'h97;
	15'h6072: q<=8'hd1;
	15'h6073: q<=8'hbd;
	15'h6074: q<=8'hd1;
	15'h6075: q<=8'hf0;
	15'h6076: q<=8'hd1;
	15'h6077: q<=8'h17;
	15'h6078: q<=8'hd2;
	15'h6079: q<=8'h75;
	15'h607a: q<=8'hd2;
	15'h607b: q<=8'he0;
	15'h607c: q<=8'hd2;
	15'h607d: q<=8'h3f;
	15'h607e: q<=8'hd3;
	15'h607f: q<=8'h79;
	15'h6080: q<=8'hd3;
	15'h6081: q<=8'hbe;
	15'h6082: q<=8'hd3;
	15'h6083: q<=8'he6;
	15'h6084: q<=8'hd3;
	15'h6085: q<=8'hff;
	15'h6086: q<=8'hd3;
	15'h6087: q<=8'h17;
	15'h6088: q<=8'hd4;
	15'h6089: q<=8'h22;
	15'h608a: q<=8'hd4;
	15'h608b: q<=8'h3a;
	15'h608c: q<=8'hd4;
	15'h608d: q<=8'h51;
	15'h608e: q<=8'hd4;
	15'h608f: q<=8'h6d;
	15'h6090: q<=8'hd4;
	15'h6091: q<=8'ha1;
	15'h6092: q<=8'hd4;
	15'h6093: q<=8'hba;
	15'h6094: q<=8'hd4;
	15'h6095: q<=8'hfd;
	15'h6096: q<=8'hd4;
	15'h6097: q<=8'h3f;
	15'h6098: q<=8'hd5;
	15'h6099: q<=8'h75;
	15'h609a: q<=8'hd5;
	15'h609b: q<=8'h85;
	15'h609c: q<=8'hd5;
	15'h609d: q<=8'ha1;
	15'h609e: q<=8'hd5;
	15'h609f: q<=8'hb9;
	15'h60a0: q<=8'hd5;
	15'h60a1: q<=8'hf6;
	15'h60a2: q<=8'hd5;
	15'h60a3: q<=8'h29;
	15'h60a4: q<=8'hd6;
	15'h60a5: q<=8'h68;
	15'h60a6: q<=8'hd6;
	15'h60a7: q<=8'h7a;
	15'h60a8: q<=8'hd6;
	15'h60a9: q<=8'h75;
	15'h60aa: q<=8'hd1;
	15'h60ab: q<=8'h9f;
	15'h60ac: q<=8'hd1;
	15'h60ad: q<=8'h9f;
	15'h60ae: q<=8'hd1;
	15'h60af: q<=8'hcf;
	15'h60b0: q<=8'hd1;
	15'h60b1: q<=8'hf6;
	15'h60b2: q<=8'hd1;
	15'h60b3: q<=8'h30;
	15'h60b4: q<=8'hd2;
	15'h60b5: q<=8'h94;
	15'h60b6: q<=8'hd2;
	15'h60b7: q<=8'hfb;
	15'h60b8: q<=8'hd2;
	15'h60b9: q<=8'h50;
	15'h60ba: q<=8'hd3;
	15'h60bb: q<=8'h8b;
	15'h60bc: q<=8'hd3;
	15'h60bd: q<=8'hcb;
	15'h60be: q<=8'hd3;
	15'h60bf: q<=8'hf5;
	15'h60c0: q<=8'hd3;
	15'h60c1: q<=8'h0e;
	15'h60c2: q<=8'hd4;
	15'h60c3: q<=8'h17;
	15'h60c4: q<=8'hd4;
	15'h60c5: q<=8'h28;
	15'h60c6: q<=8'hd4;
	15'h60c7: q<=8'h41;
	15'h60c8: q<=8'hd4;
	15'h60c9: q<=8'h5b;
	15'h60ca: q<=8'hd4;
	15'h60cb: q<=8'h83;
	15'h60cc: q<=8'hd4;
	15'h60cd: q<=8'ha1;
	15'h60ce: q<=8'hd4;
	15'h60cf: q<=8'hcc;
	15'h60d0: q<=8'hd4;
	15'h60d1: q<=8'h0e;
	15'h60d2: q<=8'hd5;
	15'h60d3: q<=8'h51;
	15'h60d4: q<=8'hd5;
	15'h60d5: q<=8'h75;
	15'h60d6: q<=8'hd5;
	15'h60d7: q<=8'h8e;
	15'h60d8: q<=8'hd5;
	15'h60d9: q<=8'ha1;
	15'h60da: q<=8'hd5;
	15'h60db: q<=8'hc8;
	15'h60dc: q<=8'hd5;
	15'h60dd: q<=8'h04;
	15'h60de: q<=8'hd6;
	15'h60df: q<=8'h3e;
	15'h60e0: q<=8'hd6;
	15'h60e1: q<=8'h6f;
	15'h60e2: q<=8'hd6;
	15'h60e3: q<=8'h8f;
	15'h60e4: q<=8'hd6;
	15'h60e5: q<=8'h7f;
	15'h60e6: q<=8'hd1;
	15'h60e7: q<=8'ha8;
	15'h60e8: q<=8'hd1;
	15'h60e9: q<=8'ha8;
	15'h60ea: q<=8'hd1;
	15'h60eb: q<=8'hde;
	15'h60ec: q<=8'hd1;
	15'h60ed: q<=8'hfc;
	15'h60ee: q<=8'hd1;
	15'h60ef: q<=8'h4d;
	15'h60f0: q<=8'hd2;
	15'h60f1: q<=8'hae;
	15'h60f2: q<=8'hd2;
	15'h60f3: q<=8'h16;
	15'h60f4: q<=8'hd3;
	15'h60f5: q<=8'h5e;
	15'h60f6: q<=8'hd3;
	15'h60f7: q<=8'ha0;
	15'h60f8: q<=8'hd3;
	15'h60f9: q<=8'hda;
	15'h60fa: q<=8'hd3;
	15'h60fb: q<=8'hed;
	15'h60fc: q<=8'hd3;
	15'h60fd: q<=8'h06;
	15'h60fe: q<=8'hd4;
	15'h60ff: q<=8'h17;
	15'h6100: q<=8'hd4;
	15'h6101: q<=8'h2d;
	15'h6102: q<=8'hd4;
	15'h6103: q<=8'h46;
	15'h6104: q<=8'hd4;
	15'h6105: q<=8'h56;
	15'h6106: q<=8'hd4;
	15'h6107: q<=8'h92;
	15'h6108: q<=8'hd4;
	15'h6109: q<=8'ha1;
	15'h610a: q<=8'hd4;
	15'h610b: q<=8'hdd;
	15'h610c: q<=8'hd4;
	15'h610d: q<=8'h1f;
	15'h610e: q<=8'hd5;
	15'h610f: q<=8'h63;
	15'h6110: q<=8'hd5;
	15'h6111: q<=8'h75;
	15'h6112: q<=8'hd5;
	15'h6113: q<=8'h97;
	15'h6114: q<=8'hd5;
	15'h6115: q<=8'ha1;
	15'h6116: q<=8'hd5;
	15'h6117: q<=8'hd9;
	15'h6118: q<=8'hd5;
	15'h6119: q<=8'h10;
	15'h611a: q<=8'hd6;
	15'h611b: q<=8'h51;
	15'h611c: q<=8'hd6;
	15'h611d: q<=8'h74;
	15'h611e: q<=8'hd6;
	15'h611f: q<=8'ha1;
	15'h6120: q<=8'hd6;
	15'h6121: q<=8'h51;
	15'h6122: q<=8'h56;
	15'h6123: q<=8'h00;
	15'h6124: q<=8'h1a;
	15'h6125: q<=8'h01;
	15'h6126: q<=8'h20;
	15'h6127: q<=8'h31;
	15'h6128: q<=8'h56;
	15'h6129: q<=8'h01;
	15'h612a: q<=8'h38;
	15'h612b: q<=8'h31;
	15'h612c: q<=8'hb0;
	15'h612d: q<=8'h41;
	15'h612e: q<=8'h00;
	15'h612f: q<=8'h11;
	15'h6130: q<=8'hf6;
	15'h6131: q<=8'h30;
	15'h6132: q<=8'h38;
	15'h6133: q<=8'h31;
	15'h6134: q<=8'hce;
	15'h6135: q<=8'h51;
	15'h6136: q<=8'h0a;
	15'h6137: q<=8'h31;
	15'h6138: q<=8'he2;
	15'h6139: q<=8'h31;
	15'h613a: q<=8'he2;
	15'h613b: q<=8'h51;
	15'h613c: q<=8'hba;
	15'h613d: q<=8'h51;
	15'h613e: q<=8'h98;
	15'h613f: q<=8'h51;
	15'h6140: q<=8'hd8;
	15'h6141: q<=8'h51;
	15'h6142: q<=8'hc9;
	15'h6143: q<=8'h31;
	15'h6144: q<=8'h56;
	15'h6145: q<=8'h51;
	15'h6146: q<=8'h80;
	15'h6147: q<=8'h51;
	15'h6148: q<=8'h80;
	15'h6149: q<=8'h51;
	15'h614a: q<=8'h80;
	15'h614b: q<=8'h51;
	15'h614c: q<=8'h80;
	15'h614d: q<=8'h71;
	15'h614e: q<=8'h92;
	15'h614f: q<=8'h51;
	15'h6150: q<=8'h80;
	15'h6151: q<=8'h31;
	15'h6152: q<=8'hb0;
	15'h6153: q<=8'h51;
	15'h6154: q<=8'h89;
	15'h6155: q<=8'h41;
	15'h6156: q<=8'h89;
	15'h6157: q<=8'h00;
	15'h6158: q<=8'h00;
	15'h6159: q<=8'h71;
	15'h615a: q<=8'h5a;
	15'h615b: q<=8'h71;
	15'h615c: q<=8'ha0;
	15'h615d: q<=8'he5;
	15'h615e: q<=8'h22;
	15'h615f: q<=8'h16;
	15'h6160: q<=8'h2e;
	15'h6161: q<=8'h1e;
	15'h6162: q<=8'h00;
	15'h6163: q<=8'h32;
	15'h6164: q<=8'h40;
	15'h6165: q<=8'h1e;
	15'h6166: q<=8'hb8;
	15'h6167: q<=8'hd9;
	15'h6168: q<=8'h20;
	15'h6169: q<=8'h26;
	15'h616a: q<=8'h30;
	15'h616b: q<=8'h00;
	15'h616c: q<=8'h1c;
	15'h616d: q<=8'h1e;
	15'h616e: q<=8'h00;
	15'h616f: q<=8'h34;
	15'h6170: q<=8'h16;
	15'h6171: q<=8'h38;
	15'h6172: q<=8'h3c;
	15'h6173: q<=8'h26;
	15'h6174: q<=8'h9e;
	15'h6175: q<=8'he5;
	15'h6176: q<=8'h3a;
	15'h6177: q<=8'h34;
	15'h6178: q<=8'h26;
	15'h6179: q<=8'h1e;
	15'h617a: q<=8'h2c;
	15'h617b: q<=8'h1e;
	15'h617c: q<=8'h30;
	15'h617d: q<=8'h1c;
	15'h617e: q<=8'h9e;
	15'h617f: q<=8'hd3;
	15'h6180: q<=8'h28;
	15'h6181: q<=8'h3e;
	15'h6182: q<=8'h1e;
	15'h6183: q<=8'h22;
	15'h6184: q<=8'h32;
	15'h6185: q<=8'h00;
	15'h6186: q<=8'h3c;
	15'h6187: q<=8'h1e;
	15'h6188: q<=8'h38;
	15'h6189: q<=8'h2e;
	15'h618a: q<=8'h26;
	15'h618b: q<=8'h30;
	15'h618c: q<=8'h16;
	15'h618d: q<=8'h1c;
	15'h618e: q<=8'hb2;
	15'h618f: q<=8'hcd;
	15'h6190: q<=8'h34;
	15'h6191: q<=8'h2c;
	15'h6192: q<=8'h16;
	15'h6193: q<=8'h46;
	15'h6194: q<=8'h1e;
	15'h6195: q<=8'h38;
	15'h6196: q<=8'h80;
	15'h6197: q<=8'hc6;
	15'h6198: q<=8'h28;
	15'h6199: q<=8'h32;
	15'h619a: q<=8'h3e;
	15'h619b: q<=8'h1e;
	15'h619c: q<=8'h3e;
	15'h619d: q<=8'h38;
	15'h619e: q<=8'h80;
	15'h619f: q<=8'hc6;
	15'h61a0: q<=8'h3a;
	15'h61a1: q<=8'h34;
	15'h61a2: q<=8'h26;
	15'h61a3: q<=8'h1e;
	15'h61a4: q<=8'h2c;
	15'h61a5: q<=8'h1e;
	15'h61a6: q<=8'h38;
	15'h61a7: q<=8'h80;
	15'h61a8: q<=8'hc6;
	15'h61a9: q<=8'h28;
	15'h61aa: q<=8'h3e;
	15'h61ab: q<=8'h22;
	15'h61ac: q<=8'h16;
	15'h61ad: q<=8'h1c;
	15'h61ae: q<=8'h32;
	15'h61af: q<=8'h38;
	15'h61b0: q<=8'h80;
	15'h61b1: q<=8'hdf;
	15'h61b2: q<=8'h34;
	15'h61b3: q<=8'h38;
	15'h61b4: q<=8'h1e;
	15'h61b5: q<=8'h3a;
	15'h61b6: q<=8'h3a;
	15'h61b7: q<=8'h00;
	15'h61b8: q<=8'h3a;
	15'h61b9: q<=8'h3c;
	15'h61ba: q<=8'h16;
	15'h61bb: q<=8'h38;
	15'h61bc: q<=8'hbc;
	15'h61bd: q<=8'hcd;
	15'h61be: q<=8'h16;
	15'h61bf: q<=8'h34;
	15'h61c0: q<=8'h34;
	15'h61c1: q<=8'h3e;
	15'h61c2: q<=8'h46;
	15'h61c3: q<=8'h1e;
	15'h61c4: q<=8'h48;
	15'h61c5: q<=8'h00;
	15'h61c6: q<=8'h3a;
	15'h61c7: q<=8'h3e;
	15'h61c8: q<=8'h38;
	15'h61c9: q<=8'h00;
	15'h61ca: q<=8'h3a;
	15'h61cb: q<=8'h3c;
	15'h61cc: q<=8'h16;
	15'h61cd: q<=8'h38;
	15'h61ce: q<=8'hbc;
	15'h61cf: q<=8'hd6;
	15'h61d0: q<=8'h3a;
	15'h61d1: q<=8'h3c;
	15'h61d2: q<=8'h16;
	15'h61d3: q<=8'h38;
	15'h61d4: q<=8'h3c;
	15'h61d5: q<=8'h00;
	15'h61d6: q<=8'h1c;
	15'h61d7: q<=8'h38;
	15'h61d8: q<=8'h3e;
	15'h61d9: q<=8'h1e;
	15'h61da: q<=8'h1a;
	15'h61db: q<=8'h2a;
	15'h61dc: q<=8'h1e;
	15'h61dd: q<=8'hb0;
	15'h61de: q<=8'hdc;
	15'h61df: q<=8'h34;
	15'h61e0: q<=8'h3e;
	15'h61e1: q<=8'h2c;
	15'h61e2: q<=8'h3a;
	15'h61e3: q<=8'h16;
	15'h61e4: q<=8'h38;
	15'h61e5: q<=8'h00;
	15'h61e6: q<=8'h3a;
	15'h61e7: q<=8'h3c;
	15'h61e8: q<=8'h16;
	15'h61e9: q<=8'h38;
	15'h61ea: q<=8'hbc;
	15'h61eb: q<=8'hf4;
	15'h61ec: q<=8'h34;
	15'h61ed: q<=8'h2c;
	15'h61ee: q<=8'h16;
	15'h61ef: q<=8'hc6;
	15'h61f0: q<=8'hf1;
	15'h61f1: q<=8'h28;
	15'h61f2: q<=8'h32;
	15'h61f3: q<=8'h3e;
	15'h61f4: q<=8'h1e;
	15'h61f5: q<=8'hc8;
	15'h61f6: q<=8'hf1;
	15'h61f7: q<=8'h3a;
	15'h61f8: q<=8'h34;
	15'h61f9: q<=8'h26;
	15'h61fa: q<=8'h1e;
	15'h61fb: q<=8'hac;
	15'h61fc: q<=8'hee;
	15'h61fd: q<=8'h28;
	15'h61fe: q<=8'h3e;
	15'h61ff: q<=8'h1e;
	15'h6200: q<=8'h22;
	15'h6201: q<=8'h3e;
	15'h6202: q<=8'h9e;
	15'h6203: q<=8'hc7;
	15'h6204: q<=8'h1e;
	15'h6205: q<=8'h30;
	15'h6206: q<=8'h3c;
	15'h6207: q<=8'h1e;
	15'h6208: q<=8'h38;
	15'h6209: q<=8'h00;
	15'h620a: q<=8'h46;
	15'h620b: q<=8'h32;
	15'h620c: q<=8'h3e;
	15'h620d: q<=8'h38;
	15'h620e: q<=8'h00;
	15'h620f: q<=8'h26;
	15'h6210: q<=8'h30;
	15'h6211: q<=8'h26;
	15'h6212: q<=8'h3c;
	15'h6213: q<=8'h26;
	15'h6214: q<=8'h16;
	15'h6215: q<=8'h2c;
	15'h6216: q<=8'hba;
	15'h6217: q<=8'hb8;
	15'h6218: q<=8'h3a;
	15'h6219: q<=8'h40;
	15'h621a: q<=8'h34;
	15'h621b: q<=8'h00;
	15'h621c: q<=8'h1e;
	15'h621d: q<=8'h30;
	15'h621e: q<=8'h3c;
	15'h621f: q<=8'h38;
	15'h6220: q<=8'h1e;
	15'h6221: q<=8'h48;
	15'h6222: q<=8'h00;
	15'h6223: q<=8'h40;
	15'h6224: q<=8'h32;
	15'h6225: q<=8'h3a;
	15'h6226: q<=8'h00;
	15'h6227: q<=8'h26;
	15'h6228: q<=8'h30;
	15'h6229: q<=8'h26;
	15'h622a: q<=8'h3c;
	15'h622b: q<=8'h26;
	15'h622c: q<=8'h16;
	15'h622d: q<=8'h2c;
	15'h622e: q<=8'h1e;
	15'h622f: q<=8'hba;
	15'h6230: q<=8'hac;
	15'h6231: q<=8'h22;
	15'h6232: q<=8'h1e;
	15'h6233: q<=8'h18;
	15'h6234: q<=8'h1e;
	15'h6235: q<=8'h30;
	15'h6236: q<=8'h00;
	15'h6237: q<=8'h3a;
	15'h6238: q<=8'h26;
	15'h6239: q<=8'h1e;
	15'h623a: q<=8'h00;
	15'h623b: q<=8'h26;
	15'h623c: q<=8'h24;
	15'h623d: q<=8'h38;
	15'h623e: q<=8'h1e;
	15'h623f: q<=8'h00;
	15'h6240: q<=8'h26;
	15'h6241: q<=8'h30;
	15'h6242: q<=8'h26;
	15'h6243: q<=8'h3c;
	15'h6244: q<=8'h26;
	15'h6245: q<=8'h16;
	15'h6246: q<=8'h2c;
	15'h6247: q<=8'h1e;
	15'h6248: q<=8'h30;
	15'h6249: q<=8'h00;
	15'h624a: q<=8'h1e;
	15'h624b: q<=8'h26;
	15'h624c: q<=8'hb0;
	15'h624d: q<=8'hc7;
	15'h624e: q<=8'h1e;
	15'h624f: q<=8'h30;
	15'h6250: q<=8'h3c;
	15'h6251: q<=8'h38;
	15'h6252: q<=8'h1e;
	15'h6253: q<=8'h00;
	15'h6254: q<=8'h3a;
	15'h6255: q<=8'h3e;
	15'h6256: q<=8'h3a;
	15'h6257: q<=8'h00;
	15'h6258: q<=8'h26;
	15'h6259: q<=8'h30;
	15'h625a: q<=8'h26;
	15'h625b: q<=8'h1a;
	15'h625c: q<=8'h26;
	15'h625d: q<=8'h16;
	15'h625e: q<=8'h2c;
	15'h625f: q<=8'h1e;
	15'h6260: q<=8'hba;
	15'h6261: q<=8'hc7;
	15'h6262: q<=8'h3a;
	15'h6263: q<=8'h34;
	15'h6264: q<=8'h26;
	15'h6265: q<=8'h30;
	15'h6266: q<=8'h00;
	15'h6267: q<=8'h2a;
	15'h6268: q<=8'h30;
	15'h6269: q<=8'h32;
	15'h626a: q<=8'h18;
	15'h626b: q<=8'h00;
	15'h626c: q<=8'h3c;
	15'h626d: q<=8'h32;
	15'h626e: q<=8'h00;
	15'h626f: q<=8'h1a;
	15'h6270: q<=8'h24;
	15'h6271: q<=8'h16;
	15'h6272: q<=8'h30;
	15'h6273: q<=8'h22;
	15'h6274: q<=8'h9e;
	15'h6275: q<=8'ha6;
	15'h6276: q<=8'h3c;
	15'h6277: q<=8'h32;
	15'h6278: q<=8'h3e;
	15'h6279: q<=8'h38;
	15'h627a: q<=8'h30;
	15'h627b: q<=8'h1e;
	15'h627c: q<=8'h48;
	15'h627d: q<=8'h00;
	15'h627e: q<=8'h2c;
	15'h627f: q<=8'h1e;
	15'h6280: q<=8'h00;
	15'h6281: q<=8'h18;
	15'h6282: q<=8'h32;
	15'h6283: q<=8'h3e;
	15'h6284: q<=8'h3c;
	15'h6285: q<=8'h32;
	15'h6286: q<=8'h30;
	15'h6287: q<=8'h00;
	15'h6288: q<=8'h34;
	15'h6289: q<=8'h32;
	15'h628a: q<=8'h3e;
	15'h628b: q<=8'h38;
	15'h628c: q<=8'h00;
	15'h628d: q<=8'h1a;
	15'h628e: q<=8'h24;
	15'h628f: q<=8'h16;
	15'h6290: q<=8'h30;
	15'h6291: q<=8'h22;
	15'h6292: q<=8'h1e;
	15'h6293: q<=8'hb8;
	15'h6294: q<=8'hb5;
	15'h6295: q<=8'h2a;
	15'h6296: q<=8'h30;
	15'h6297: q<=8'h32;
	15'h6298: q<=8'h34;
	15'h6299: q<=8'h20;
	15'h629a: q<=8'h00;
	15'h629b: q<=8'h1c;
	15'h629c: q<=8'h38;
	15'h629d: q<=8'h1e;
	15'h629e: q<=8'h24;
	15'h629f: q<=8'h1e;
	15'h62a0: q<=8'h30;
	15'h62a1: q<=8'h00;
	15'h62a2: q<=8'h48;
	15'h62a3: q<=8'h3e;
	15'h62a4: q<=8'h2e;
	15'h62a5: q<=8'h00;
	15'h62a6: q<=8'h42;
	15'h62a7: q<=8'h1e;
	15'h62a8: q<=8'h1a;
	15'h62a9: q<=8'h24;
	15'h62aa: q<=8'h3a;
	15'h62ab: q<=8'h1e;
	15'h62ac: q<=8'h2c;
	15'h62ad: q<=8'hb0;
	15'h62ae: q<=8'hac;
	15'h62af: q<=8'h22;
	15'h62b0: q<=8'h26;
	15'h62b1: q<=8'h38;
	15'h62b2: q<=8'h1e;
	15'h62b3: q<=8'h00;
	15'h62b4: q<=8'h2c;
	15'h62b5: q<=8'h16;
	15'h62b6: q<=8'h00;
	15'h62b7: q<=8'h34;
	15'h62b8: q<=8'h1e;
	15'h62b9: q<=8'h38;
	15'h62ba: q<=8'h26;
	15'h62bb: q<=8'h2c;
	15'h62bc: q<=8'h2c;
	15'h62bd: q<=8'h16;
	15'h62be: q<=8'h00;
	15'h62bf: q<=8'h34;
	15'h62c0: q<=8'h16;
	15'h62c1: q<=8'h38;
	15'h62c2: q<=8'h16;
	15'h62c3: q<=8'h00;
	15'h62c4: q<=8'h1a;
	15'h62c5: q<=8'h16;
	15'h62c6: q<=8'h2e;
	15'h62c7: q<=8'h18;
	15'h62c8: q<=8'h26;
	15'h62c9: q<=8'h16;
	15'h62ca: q<=8'hb8;
	15'h62cb: q<=8'hc4;
	15'h62cc: q<=8'h34;
	15'h62cd: q<=8'h38;
	15'h62ce: q<=8'h1e;
	15'h62cf: q<=8'h3a;
	15'h62d0: q<=8'h3a;
	15'h62d1: q<=8'h00;
	15'h62d2: q<=8'h20;
	15'h62d3: q<=8'h26;
	15'h62d4: q<=8'h38;
	15'h62d5: q<=8'h1e;
	15'h62d6: q<=8'h00;
	15'h62d7: q<=8'h3c;
	15'h62d8: q<=8'h32;
	15'h62d9: q<=8'h00;
	15'h62da: q<=8'h3a;
	15'h62db: q<=8'h1e;
	15'h62dc: q<=8'h2c;
	15'h62dd: q<=8'h1e;
	15'h62de: q<=8'h1a;
	15'h62df: q<=8'hbc;
	15'h62e0: q<=8'hb2;
	15'h62e1: q<=8'h34;
	15'h62e2: q<=8'h32;
	15'h62e3: q<=8'h3e;
	15'h62e4: q<=8'h3a;
	15'h62e5: q<=8'h3a;
	15'h62e6: q<=8'h1e;
	15'h62e7: q<=8'h48;
	15'h62e8: q<=8'h00;
	15'h62e9: q<=8'h20;
	15'h62ea: q<=8'h1e;
	15'h62eb: q<=8'h3e;
	15'h62ec: q<=8'h00;
	15'h62ed: q<=8'h36;
	15'h62ee: q<=8'h3e;
	15'h62ef: q<=8'h16;
	15'h62f0: q<=8'h30;
	15'h62f1: q<=8'h1c;
	15'h62f2: q<=8'h00;
	15'h62f3: q<=8'h1a;
	15'h62f4: q<=8'h32;
	15'h62f5: q<=8'h38;
	15'h62f6: q<=8'h38;
	15'h62f7: q<=8'h1e;
	15'h62f8: q<=8'h1a;
	15'h62f9: q<=8'h3c;
	15'h62fa: q<=8'h9e;
	15'h62fb: q<=8'hb2;
	15'h62fc: q<=8'h20;
	15'h62fd: q<=8'h26;
	15'h62fe: q<=8'h38;
	15'h62ff: q<=8'h1e;
	15'h6300: q<=8'h00;
	15'h6301: q<=8'h1c;
	15'h6302: q<=8'h38;
	15'h6303: q<=8'h3e;
	15'h6304: q<=8'h1e;
	15'h6305: q<=8'h1a;
	15'h6306: q<=8'h2a;
	15'h6307: q<=8'h1e;
	15'h6308: q<=8'h30;
	15'h6309: q<=8'h00;
	15'h630a: q<=8'h42;
	15'h630b: q<=8'h1e;
	15'h630c: q<=8'h30;
	15'h630d: q<=8'h30;
	15'h630e: q<=8'h00;
	15'h630f: q<=8'h38;
	15'h6310: q<=8'h26;
	15'h6311: q<=8'h1a;
	15'h6312: q<=8'h24;
	15'h6313: q<=8'h3c;
	15'h6314: q<=8'h26;
	15'h6315: q<=8'ha2;
	15'h6316: q<=8'hac;
	15'h6317: q<=8'h32;
	15'h6318: q<=8'h34;
	15'h6319: q<=8'h38;
	15'h631a: q<=8'h26;
	15'h631b: q<=8'h2e;
	15'h631c: q<=8'h16;
	15'h631d: q<=8'h00;
	15'h631e: q<=8'h20;
	15'h631f: q<=8'h26;
	15'h6320: q<=8'h38;
	15'h6321: q<=8'h1e;
	15'h6322: q<=8'h00;
	15'h6323: q<=8'h34;
	15'h6324: q<=8'h16;
	15'h6325: q<=8'h38;
	15'h6326: q<=8'h16;
	15'h6327: q<=8'h00;
	15'h6328: q<=8'h3a;
	15'h6329: q<=8'h1e;
	15'h632a: q<=8'h2c;
	15'h632b: q<=8'h1e;
	15'h632c: q<=8'h1a;
	15'h632d: q<=8'h1a;
	15'h632e: q<=8'h26;
	15'h632f: q<=8'h32;
	15'h6330: q<=8'h30;
	15'h6331: q<=8'h16;
	15'h6332: q<=8'hb8;
	15'h6333: q<=8'hbc;
	15'h6334: q<=8'h24;
	15'h6335: q<=8'h26;
	15'h6336: q<=8'h22;
	15'h6337: q<=8'h24;
	15'h6338: q<=8'h00;
	15'h6339: q<=8'h3a;
	15'h633a: q<=8'h1a;
	15'h633b: q<=8'h32;
	15'h633c: q<=8'h38;
	15'h633d: q<=8'h1e;
	15'h633e: q<=8'hba;
	15'h633f: q<=8'h9e;
	15'h6340: q<=8'h2e;
	15'h6341: q<=8'h1e;
	15'h6342: q<=8'h26;
	15'h6343: q<=8'h2c;
	15'h6344: q<=8'h2c;
	15'h6345: q<=8'h1e;
	15'h6346: q<=8'h3e;
	15'h6347: q<=8'h38;
	15'h6348: q<=8'h3a;
	15'h6349: q<=8'h00;
	15'h634a: q<=8'h3a;
	15'h634b: q<=8'h1a;
	15'h634c: q<=8'h32;
	15'h634d: q<=8'h38;
	15'h634e: q<=8'h1e;
	15'h634f: q<=8'hba;
	15'h6350: q<=8'hb0;
	15'h6351: q<=8'h24;
	15'h6352: q<=8'h32;
	15'h6353: q<=8'h1e;
	15'h6354: q<=8'h1a;
	15'h6355: q<=8'h24;
	15'h6356: q<=8'h3a;
	15'h6357: q<=8'h3c;
	15'h6358: q<=8'h48;
	15'h6359: q<=8'h16;
	15'h635a: q<=8'h24;
	15'h635b: q<=8'h2c;
	15'h635c: q<=8'h1e;
	15'h635d: q<=8'hb0;
	15'h635e: q<=8'hd4;
	15'h635f: q<=8'h38;
	15'h6360: q<=8'h1e;
	15'h6361: q<=8'h1a;
	15'h6362: q<=8'h32;
	15'h6363: q<=8'h38;
	15'h6364: q<=8'h1c;
	15'h6365: q<=8'hba;
	15'h6366: q<=8'hc2;
	15'h6367: q<=8'h38;
	15'h6368: q<=8'h16;
	15'h6369: q<=8'h30;
	15'h636a: q<=8'h2a;
	15'h636b: q<=8'h26;
	15'h636c: q<=8'h30;
	15'h636d: q<=8'h22;
	15'h636e: q<=8'h00;
	15'h636f: q<=8'h20;
	15'h6370: q<=8'h38;
	15'h6371: q<=8'h32;
	15'h6372: q<=8'h2e;
	15'h6373: q<=8'h00;
	15'h6374: q<=8'h04;
	15'h6375: q<=8'h00;
	15'h6376: q<=8'h3c;
	15'h6377: q<=8'h32;
	15'h6378: q<=8'h80;
	15'h6379: q<=8'hc2;
	15'h637a: q<=8'h34;
	15'h637b: q<=8'h2c;
	15'h637c: q<=8'h16;
	15'h637d: q<=8'h1a;
	15'h637e: q<=8'h1e;
	15'h637f: q<=8'h2e;
	15'h6380: q<=8'h1e;
	15'h6381: q<=8'h30;
	15'h6382: q<=8'h3c;
	15'h6383: q<=8'h00;
	15'h6384: q<=8'h1c;
	15'h6385: q<=8'h1e;
	15'h6386: q<=8'h00;
	15'h6387: q<=8'h04;
	15'h6388: q<=8'h00;
	15'h6389: q<=8'h16;
	15'h638a: q<=8'h80;
	15'h638b: q<=8'hbc;
	15'h638c: q<=8'h38;
	15'h638d: q<=8'h16;
	15'h638e: q<=8'h30;
	15'h638f: q<=8'h22;
	15'h6390: q<=8'h2c;
	15'h6391: q<=8'h26;
	15'h6392: q<=8'h3a;
	15'h6393: q<=8'h3c;
	15'h6394: q<=8'h1e;
	15'h6395: q<=8'h00;
	15'h6396: q<=8'h40;
	15'h6397: q<=8'h32;
	15'h6398: q<=8'h30;
	15'h6399: q<=8'h00;
	15'h639a: q<=8'h04;
	15'h639b: q<=8'h00;
	15'h639c: q<=8'h48;
	15'h639d: q<=8'h3e;
	15'h639e: q<=8'h2e;
	15'h639f: q<=8'h80;
	15'h63a0: q<=8'hc8;
	15'h63a1: q<=8'h38;
	15'h63a2: q<=8'h16;
	15'h63a3: q<=8'h30;
	15'h63a4: q<=8'h2a;
	15'h63a5: q<=8'h26;
	15'h63a6: q<=8'h30;
	15'h63a7: q<=8'h22;
	15'h63a8: q<=8'h00;
	15'h63a9: q<=8'h1c;
	15'h63aa: q<=8'h1e;
	15'h63ab: q<=8'h00;
	15'h63ac: q<=8'h04;
	15'h63ad: q<=8'h00;
	15'h63ae: q<=8'h16;
	15'h63af: q<=8'h80;
	15'h63b0: q<=8'hd9;
	15'h63b1: q<=8'h38;
	15'h63b2: q<=8'h16;
	15'h63b3: q<=8'h3c;
	15'h63b4: q<=8'h1e;
	15'h63b5: q<=8'h00;
	15'h63b6: q<=8'h46;
	15'h63b7: q<=8'h32;
	15'h63b8: q<=8'h3e;
	15'h63b9: q<=8'h38;
	15'h63ba: q<=8'h3a;
	15'h63bb: q<=8'h1e;
	15'h63bc: q<=8'h2c;
	15'h63bd: q<=8'ha0;
	15'h63be: q<=8'hdc;
	15'h63bf: q<=8'h1e;
	15'h63c0: q<=8'h40;
	15'h63c1: q<=8'h16;
	15'h63c2: q<=8'h2c;
	15'h63c3: q<=8'h3e;
	15'h63c4: q<=8'h1e;
	15'h63c5: q<=8'h48;
	15'h63c6: q<=8'h4c;
	15'h63c7: q<=8'h40;
	15'h63c8: q<=8'h32;
	15'h63c9: q<=8'h3e;
	15'h63ca: q<=8'hba;
	15'h63cb: q<=8'hd6;
	15'h63cc: q<=8'h3a;
	15'h63cd: q<=8'h1e;
	15'h63ce: q<=8'h2c;
	15'h63cf: q<=8'h18;
	15'h63d0: q<=8'h3a;
	15'h63d1: q<=8'h3c;
	15'h63d2: q<=8'h00;
	15'h63d3: q<=8'h38;
	15'h63d4: q<=8'h1e;
	15'h63d5: q<=8'h1a;
	15'h63d6: q<=8'h24;
	15'h63d7: q<=8'h30;
	15'h63d8: q<=8'h1e;
	15'h63d9: q<=8'hb0;
	15'h63da: q<=8'hdf;
	15'h63db: q<=8'h1a;
	15'h63dc: q<=8'h16;
	15'h63dd: q<=8'h2c;
	15'h63de: q<=8'h26;
	15'h63df: q<=8'h20;
	15'h63e0: q<=8'h26;
	15'h63e1: q<=8'h36;
	15'h63e2: q<=8'h3e;
	15'h63e3: q<=8'h1e;
	15'h63e4: q<=8'h3a;
	15'h63e5: q<=8'h9e;
	15'h63e6: q<=8'haa;
	15'h63e7: q<=8'h30;
	15'h63e8: q<=8'h32;
	15'h63e9: q<=8'h40;
	15'h63ea: q<=8'h26;
	15'h63eb: q<=8'h1a;
	15'h63ec: q<=8'h9e;
	15'h63ed: q<=8'haa;
	15'h63ee: q<=8'h30;
	15'h63ef: q<=8'h32;
	15'h63f0: q<=8'h40;
	15'h63f1: q<=8'h26;
	15'h63f2: q<=8'h1a;
	15'h63f3: q<=8'h26;
	15'h63f4: q<=8'hb2;
	15'h63f5: q<=8'haa;
	15'h63f6: q<=8'h16;
	15'h63f7: q<=8'h30;
	15'h63f8: q<=8'h20;
	15'h63f9: q<=8'h16;
	15'h63fa: q<=8'h1e;
	15'h63fb: q<=8'h30;
	15'h63fc: q<=8'h22;
	15'h63fd: q<=8'h1e;
	15'h63fe: q<=8'hb8;
	15'h63ff: q<=8'h4a;
	15'h6400: q<=8'h1e;
	15'h6401: q<=8'h44;
	15'h6402: q<=8'h34;
	15'h6403: q<=8'h1e;
	15'h6404: q<=8'h38;
	15'h6405: q<=8'hbc;
	15'h6406: q<=8'h45;
	15'h6407: q<=8'h1e;
	15'h6408: q<=8'h44;
	15'h6409: q<=8'h34;
	15'h640a: q<=8'h1e;
	15'h640b: q<=8'h38;
	15'h640c: q<=8'h3c;
	15'h640d: q<=8'hb2;
	15'h640e: q<=8'h40;
	15'h640f: q<=8'h1e;
	15'h6410: q<=8'h38;
	15'h6411: q<=8'h20;
	15'h6412: q<=8'h16;
	15'h6413: q<=8'h24;
	15'h6414: q<=8'h38;
	15'h6415: q<=8'h1e;
	15'h6416: q<=8'hb0;
	15'h6417: q<=8'h8b;
	15'h6418: q<=8'h18;
	15'h6419: q<=8'h32;
	15'h641a: q<=8'h30;
	15'h641b: q<=8'h3e;
	15'h641c: q<=8'hba;
	15'h641d: q<=8'he8;
	15'h641e: q<=8'h3c;
	15'h641f: q<=8'h26;
	15'h6420: q<=8'h2e;
	15'h6421: q<=8'h9e;
	15'h6422: q<=8'he0;
	15'h6423: q<=8'h1c;
	15'h6424: q<=8'h3e;
	15'h6425: q<=8'h38;
	15'h6426: q<=8'h1e;
	15'h6427: q<=8'h9e;
	15'h6428: q<=8'he8;
	15'h6429: q<=8'h48;
	15'h642a: q<=8'h1e;
	15'h642b: q<=8'h26;
	15'h642c: q<=8'hbc;
	15'h642d: q<=8'he4;
	15'h642e: q<=8'h3c;
	15'h642f: q<=8'h26;
	15'h6430: q<=8'h1e;
	15'h6431: q<=8'h2e;
	15'h6432: q<=8'h34;
	15'h6433: q<=8'hb2;
	15'h6434: q<=8'h8b;
	15'h6435: q<=8'h2c;
	15'h6436: q<=8'h1e;
	15'h6437: q<=8'h40;
	15'h6438: q<=8'h1e;
	15'h6439: q<=8'hac;
	15'h643a: q<=8'h8b;
	15'h643b: q<=8'h30;
	15'h643c: q<=8'h26;
	15'h643d: q<=8'h40;
	15'h643e: q<=8'h1e;
	15'h643f: q<=8'h16;
	15'h6440: q<=8'hbe;
	15'h6441: q<=8'h8b;
	15'h6442: q<=8'h22;
	15'h6443: q<=8'h38;
	15'h6444: q<=8'h16;
	15'h6445: q<=8'h9c;
	15'h6446: q<=8'h8b;
	15'h6447: q<=8'h30;
	15'h6448: q<=8'h26;
	15'h6449: q<=8'h40;
	15'h644a: q<=8'h1e;
	15'h644b: q<=8'hac;
	15'h644c: q<=8'h8b;
	15'h644d: q<=8'h24;
	15'h644e: q<=8'h32;
	15'h644f: q<=8'h2c;
	15'h6450: q<=8'h9e;
	15'h6451: q<=8'h8b;
	15'h6452: q<=8'h3c;
	15'h6453: q<=8'h38;
	15'h6454: q<=8'h32;
	15'h6455: q<=8'hbe;
	15'h6456: q<=8'h8b;
	15'h6457: q<=8'h24;
	15'h6458: q<=8'h32;
	15'h6459: q<=8'h46;
	15'h645a: q<=8'hb2;
	15'h645b: q<=8'h8b;
	15'h645c: q<=8'h2c;
	15'h645d: q<=8'h32;
	15'h645e: q<=8'h1a;
	15'h645f: q<=8'ha4;
	15'h6460: q<=8'hdc;
	15'h6461: q<=8'h26;
	15'h6462: q<=8'h30;
	15'h6463: q<=8'h3a;
	15'h6464: q<=8'h1e;
	15'h6465: q<=8'h38;
	15'h6466: q<=8'h3c;
	15'h6467: q<=8'h00;
	15'h6468: q<=8'h1a;
	15'h6469: q<=8'h32;
	15'h646a: q<=8'h26;
	15'h646b: q<=8'h30;
	15'h646c: q<=8'hba;
	15'h646d: q<=8'hc1;
	15'h646e: q<=8'h26;
	15'h646f: q<=8'h30;
	15'h6470: q<=8'h3c;
	15'h6471: q<=8'h38;
	15'h6472: q<=8'h32;
	15'h6473: q<=8'h1c;
	15'h6474: q<=8'h3e;
	15'h6475: q<=8'h26;
	15'h6476: q<=8'h38;
	15'h6477: q<=8'h1e;
	15'h6478: q<=8'h00;
	15'h6479: q<=8'h2c;
	15'h647a: q<=8'h1e;
	15'h647b: q<=8'h3a;
	15'h647c: q<=8'h00;
	15'h647d: q<=8'h34;
	15'h647e: q<=8'h26;
	15'h647f: q<=8'h1e;
	15'h6480: q<=8'h1a;
	15'h6481: q<=8'h1e;
	15'h6482: q<=8'hba;
	15'h6483: q<=8'hd6;
	15'h6484: q<=8'h22;
	15'h6485: q<=8'h1e;
	15'h6486: q<=8'h2c;
	15'h6487: q<=8'h1c;
	15'h6488: q<=8'h00;
	15'h6489: q<=8'h1e;
	15'h648a: q<=8'h26;
	15'h648b: q<=8'h30;
	15'h648c: q<=8'h42;
	15'h648d: q<=8'h1e;
	15'h648e: q<=8'h38;
	15'h648f: q<=8'h20;
	15'h6490: q<=8'h1e;
	15'h6491: q<=8'hb0;
	15'h6492: q<=8'hd6;
	15'h6493: q<=8'h26;
	15'h6494: q<=8'h30;
	15'h6495: q<=8'h3a;
	15'h6496: q<=8'h1e;
	15'h6497: q<=8'h38;
	15'h6498: q<=8'h3c;
	15'h6499: q<=8'h1e;
	15'h649a: q<=8'h00;
	15'h649b: q<=8'h20;
	15'h649c: q<=8'h26;
	15'h649d: q<=8'h1a;
	15'h649e: q<=8'h24;
	15'h649f: q<=8'h16;
	15'h64a0: q<=8'hba;
	15'h64a1: q<=8'h00;
	15'h64a2: q<=8'h20;
	15'h64a3: q<=8'h38;
	15'h64a4: q<=8'h1e;
	15'h64a5: q<=8'h1e;
	15'h64a6: q<=8'h00;
	15'h64a7: q<=8'h34;
	15'h64a8: q<=8'h2c;
	15'h64a9: q<=8'h16;
	15'h64aa: q<=8'hc6;
	15'h64ab: q<=8'h0e;
	15'h64ac: q<=8'h04;
	15'h64ad: q<=8'h00;
	15'h64ae: q<=8'h1a;
	15'h64af: q<=8'h32;
	15'h64b0: q<=8'h26;
	15'h64b1: q<=8'h30;
	15'h64b2: q<=8'h00;
	15'h64b3: q<=8'h06;
	15'h64b4: q<=8'h00;
	15'h64b5: q<=8'h34;
	15'h64b6: q<=8'h2c;
	15'h64b7: q<=8'h16;
	15'h64b8: q<=8'h46;
	15'h64b9: q<=8'hba;
	15'h64ba: q<=8'hfa;
	15'h64bb: q<=8'h04;
	15'h64bc: q<=8'h00;
	15'h64bd: q<=8'h34;
	15'h64be: q<=8'h26;
	15'h64bf: q<=8'h1e;
	15'h64c0: q<=8'h1a;
	15'h64c1: q<=8'h1e;
	15'h64c2: q<=8'h00;
	15'h64c3: q<=8'h06;
	15'h64c4: q<=8'h00;
	15'h64c5: q<=8'h28;
	15'h64c6: q<=8'h32;
	15'h64c7: q<=8'h3e;
	15'h64c8: q<=8'h1e;
	15'h64c9: q<=8'h3e;
	15'h64ca: q<=8'h38;
	15'h64cb: q<=8'hba;
	15'h64cc: q<=8'h00;
	15'h64cd: q<=8'h04;
	15'h64ce: q<=8'h00;
	15'h64cf: q<=8'h2e;
	15'h64d0: q<=8'h3e;
	15'h64d1: q<=8'h1e;
	15'h64d2: q<=8'h30;
	15'h64d3: q<=8'h48;
	15'h64d4: q<=8'h00;
	15'h64d5: q<=8'h06;
	15'h64d6: q<=8'h00;
	15'h64d7: q<=8'h3a;
	15'h64d8: q<=8'h34;
	15'h64d9: q<=8'h26;
	15'h64da: q<=8'h1e;
	15'h64db: q<=8'h2c;
	15'h64dc: q<=8'h9e;
	15'h64dd: q<=8'hfa;
	15'h64de: q<=8'h04;
	15'h64df: q<=8'h00;
	15'h64e0: q<=8'h2e;
	15'h64e1: q<=8'h32;
	15'h64e2: q<=8'h30;
	15'h64e3: q<=8'h1e;
	15'h64e4: q<=8'h1c;
	15'h64e5: q<=8'h16;
	15'h64e6: q<=8'h00;
	15'h64e7: q<=8'h06;
	15'h64e8: q<=8'h00;
	15'h64e9: q<=8'h28;
	15'h64ea: q<=8'h3e;
	15'h64eb: q<=8'h1e;
	15'h64ec: q<=8'h22;
	15'h64ed: q<=8'h32;
	15'h64ee: q<=8'hba;
	15'h64ef: q<=8'h14;
	15'h64f0: q<=8'h04;
	15'h64f1: q<=8'h00;
	15'h64f2: q<=8'h1a;
	15'h64f3: q<=8'h32;
	15'h64f4: q<=8'h26;
	15'h64f5: q<=8'h30;
	15'h64f6: q<=8'h00;
	15'h64f7: q<=8'h04;
	15'h64f8: q<=8'h00;
	15'h64f9: q<=8'h34;
	15'h64fa: q<=8'h2c;
	15'h64fb: q<=8'h16;
	15'h64fc: q<=8'hc6;
	15'h64fd: q<=8'h00;
	15'h64fe: q<=8'h04;
	15'h64ff: q<=8'h00;
	15'h6500: q<=8'h34;
	15'h6501: q<=8'h26;
	15'h6502: q<=8'h1e;
	15'h6503: q<=8'h1a;
	15'h6504: q<=8'h1e;
	15'h6505: q<=8'h00;
	15'h6506: q<=8'h04;
	15'h6507: q<=8'h00;
	15'h6508: q<=8'h28;
	15'h6509: q<=8'h32;
	15'h650a: q<=8'h3e;
	15'h650b: q<=8'h1e;
	15'h650c: q<=8'h3e;
	15'h650d: q<=8'hb8;
	15'h650e: q<=8'h00;
	15'h650f: q<=8'h04;
	15'h6510: q<=8'h00;
	15'h6511: q<=8'h2e;
	15'h6512: q<=8'h3e;
	15'h6513: q<=8'h1e;
	15'h6514: q<=8'h30;
	15'h6515: q<=8'h48;
	15'h6516: q<=8'h1e;
	15'h6517: q<=8'h00;
	15'h6518: q<=8'h04;
	15'h6519: q<=8'h00;
	15'h651a: q<=8'h3a;
	15'h651b: q<=8'h34;
	15'h651c: q<=8'h26;
	15'h651d: q<=8'h1e;
	15'h651e: q<=8'hac;
	15'h651f: q<=8'h00;
	15'h6520: q<=8'h04;
	15'h6521: q<=8'h00;
	15'h6522: q<=8'h2e;
	15'h6523: q<=8'h32;
	15'h6524: q<=8'h30;
	15'h6525: q<=8'h1e;
	15'h6526: q<=8'h1c;
	15'h6527: q<=8'h16;
	15'h6528: q<=8'h00;
	15'h6529: q<=8'h04;
	15'h652a: q<=8'h00;
	15'h652b: q<=8'h28;
	15'h652c: q<=8'h3e;
	15'h652d: q<=8'h1e;
	15'h652e: q<=8'h22;
	15'h652f: q<=8'hb2;
	15'h6530: q<=8'h0e;
	15'h6531: q<=8'h06;
	15'h6532: q<=8'h00;
	15'h6533: q<=8'h1a;
	15'h6534: q<=8'h32;
	15'h6535: q<=8'h26;
	15'h6536: q<=8'h30;
	15'h6537: q<=8'h3a;
	15'h6538: q<=8'h00;
	15'h6539: q<=8'h04;
	15'h653a: q<=8'h00;
	15'h653b: q<=8'h34;
	15'h653c: q<=8'h2c;
	15'h653d: q<=8'h16;
	15'h653e: q<=8'hc6;
	15'h653f: q<=8'hfa;
	15'h6540: q<=8'h06;
	15'h6541: q<=8'h00;
	15'h6542: q<=8'h34;
	15'h6543: q<=8'h26;
	15'h6544: q<=8'h1e;
	15'h6545: q<=8'h1a;
	15'h6546: q<=8'h1e;
	15'h6547: q<=8'h3a;
	15'h6548: q<=8'h00;
	15'h6549: q<=8'h04;
	15'h654a: q<=8'h00;
	15'h654b: q<=8'h28;
	15'h654c: q<=8'h32;
	15'h654d: q<=8'h3e;
	15'h654e: q<=8'h1e;
	15'h654f: q<=8'h3e;
	15'h6550: q<=8'hb8;
	15'h6551: q<=8'hfa;
	15'h6552: q<=8'h06;
	15'h6553: q<=8'h00;
	15'h6554: q<=8'h2e;
	15'h6555: q<=8'h3e;
	15'h6556: q<=8'h1e;
	15'h6557: q<=8'h30;
	15'h6558: q<=8'h48;
	15'h6559: q<=8'h1e;
	15'h655a: q<=8'h30;
	15'h655b: q<=8'h00;
	15'h655c: q<=8'h04;
	15'h655d: q<=8'h00;
	15'h655e: q<=8'h3a;
	15'h655f: q<=8'h34;
	15'h6560: q<=8'h26;
	15'h6561: q<=8'h1e;
	15'h6562: q<=8'hac;
	15'h6563: q<=8'hfa;
	15'h6564: q<=8'h06;
	15'h6565: q<=8'h00;
	15'h6566: q<=8'h2e;
	15'h6567: q<=8'h32;
	15'h6568: q<=8'h30;
	15'h6569: q<=8'h1e;
	15'h656a: q<=8'h1c;
	15'h656b: q<=8'h16;
	15'h656c: q<=8'h3a;
	15'h656d: q<=8'h00;
	15'h656e: q<=8'h04;
	15'h656f: q<=8'h00;
	15'h6570: q<=8'h28;
	15'h6571: q<=8'h3e;
	15'h6572: q<=8'h1e;
	15'h6573: q<=8'h22;
	15'h6574: q<=8'hb2;
	15'h6575: q<=8'hd3;
	15'h6576: q<=8'h50;
	15'h6577: q<=8'h00;
	15'h6578: q<=8'h2e;
	15'h6579: q<=8'h1a;
	15'h657a: q<=8'h2e;
	15'h657b: q<=8'h2c;
	15'h657c: q<=8'h44;
	15'h657d: q<=8'h44;
	15'h657e: q<=8'h44;
	15'h657f: q<=8'h00;
	15'h6580: q<=8'h16;
	15'h6581: q<=8'h3c;
	15'h6582: q<=8'h16;
	15'h6583: q<=8'h38;
	15'h6584: q<=8'ha6;
	15'h6585: q<=8'ha0;
	15'h6586: q<=8'h1a;
	15'h6587: q<=8'h38;
	15'h6588: q<=8'h1e;
	15'h6589: q<=8'h1c;
	15'h658a: q<=8'h26;
	15'h658b: q<=8'h3c;
	15'h658c: q<=8'h3a;
	15'h658d: q<=8'h80;
	15'h658e: q<=8'ha0;
	15'h658f: q<=8'h2a;
	15'h6590: q<=8'h38;
	15'h6591: q<=8'h1e;
	15'h6592: q<=8'h1c;
	15'h6593: q<=8'h26;
	15'h6594: q<=8'h3c;
	15'h6595: q<=8'h1e;
	15'h6596: q<=8'h80;
	15'h6597: q<=8'ha0;
	15'h6598: q<=8'h1a;
	15'h6599: q<=8'h38;
	15'h659a: q<=8'h1e;
	15'h659b: q<=8'h1c;
	15'h659c: q<=8'h26;
	15'h659d: q<=8'h3c;
	15'h659e: q<=8'h32;
	15'h659f: q<=8'h3a;
	15'h65a0: q<=8'h80;
	15'h65a1: q<=8'hda;
	15'h65a2: q<=8'h18;
	15'h65a3: q<=8'h32;
	15'h65a4: q<=8'h30;
	15'h65a5: q<=8'h3e;
	15'h65a6: q<=8'h3a;
	15'h65a7: q<=8'h80;
	15'h65a8: q<=8'hd0;
	15'h65a9: q<=8'h06;
	15'h65aa: q<=8'h00;
	15'h65ab: q<=8'h1a;
	15'h65ac: q<=8'h38;
	15'h65ad: q<=8'h1e;
	15'h65ae: q<=8'h1c;
	15'h65af: q<=8'h26;
	15'h65b0: q<=8'h3c;
	15'h65b1: q<=8'h00;
	15'h65b2: q<=8'h2e;
	15'h65b3: q<=8'h26;
	15'h65b4: q<=8'h30;
	15'h65b5: q<=8'h26;
	15'h65b6: q<=8'h2e;
	15'h65b7: q<=8'h3e;
	15'h65b8: q<=8'hae;
	15'h65b9: q<=8'hd6;
	15'h65ba: q<=8'h06;
	15'h65bb: q<=8'h00;
	15'h65bc: q<=8'h28;
	15'h65bd: q<=8'h1e;
	15'h65be: q<=8'h3e;
	15'h65bf: q<=8'h44;
	15'h65c0: q<=8'h00;
	15'h65c1: q<=8'h2e;
	15'h65c2: q<=8'h26;
	15'h65c3: q<=8'h30;
	15'h65c4: q<=8'h26;
	15'h65c5: q<=8'h2e;
	15'h65c6: q<=8'h3e;
	15'h65c7: q<=8'hae;
	15'h65c8: q<=8'hd0;
	15'h65c9: q<=8'h06;
	15'h65ca: q<=8'h00;
	15'h65cb: q<=8'h3a;
	15'h65cc: q<=8'h34;
	15'h65cd: q<=8'h26;
	15'h65ce: q<=8'h1e;
	15'h65cf: q<=8'h2c;
	15'h65d0: q<=8'h1e;
	15'h65d1: q<=8'h00;
	15'h65d2: q<=8'h2e;
	15'h65d3: q<=8'h26;
	15'h65d4: q<=8'h30;
	15'h65d5: q<=8'h26;
	15'h65d6: q<=8'h2e;
	15'h65d7: q<=8'h3e;
	15'h65d8: q<=8'hae;
	15'h65d9: q<=8'hd3;
	15'h65da: q<=8'h06;
	15'h65db: q<=8'h00;
	15'h65dc: q<=8'h28;
	15'h65dd: q<=8'h3e;
	15'h65de: q<=8'h1e;
	15'h65df: q<=8'h22;
	15'h65e0: q<=8'h32;
	15'h65e1: q<=8'h3a;
	15'h65e2: q<=8'h00;
	15'h65e3: q<=8'h2e;
	15'h65e4: q<=8'h26;
	15'h65e5: q<=8'h30;
	15'h65e6: q<=8'h26;
	15'h65e7: q<=8'h2e;
	15'h65e8: q<=8'hb2;
	15'h65e9: q<=8'hc8;
	15'h65ea: q<=8'h18;
	15'h65eb: q<=8'h32;
	15'h65ec: q<=8'h30;
	15'h65ed: q<=8'h3e;
	15'h65ee: q<=8'h3a;
	15'h65ef: q<=8'h00;
	15'h65f0: q<=8'h1e;
	15'h65f1: q<=8'h40;
	15'h65f2: q<=8'h1e;
	15'h65f3: q<=8'h38;
	15'h65f4: q<=8'h46;
	15'h65f5: q<=8'h80;
	15'h65f6: q<=8'hce;
	15'h65f7: q<=8'h18;
	15'h65f8: q<=8'h32;
	15'h65f9: q<=8'h30;
	15'h65fa: q<=8'h3e;
	15'h65fb: q<=8'h3a;
	15'h65fc: q<=8'h00;
	15'h65fd: q<=8'h1a;
	15'h65fe: q<=8'h24;
	15'h65ff: q<=8'h16;
	15'h6600: q<=8'h36;
	15'h6601: q<=8'h3e;
	15'h6602: q<=8'h1e;
	15'h6603: q<=8'h80;
	15'h6604: q<=8'hce;
	15'h6605: q<=8'h18;
	15'h6606: q<=8'h32;
	15'h6607: q<=8'h30;
	15'h6608: q<=8'h3e;
	15'h6609: q<=8'h3a;
	15'h660a: q<=8'h00;
	15'h660b: q<=8'h28;
	15'h660c: q<=8'h1e;
	15'h660d: q<=8'h1c;
	15'h660e: q<=8'h1e;
	15'h660f: q<=8'h80;
	15'h6610: q<=8'hc8;
	15'h6611: q<=8'h18;
	15'h6612: q<=8'h32;
	15'h6613: q<=8'h30;
	15'h6614: q<=8'h3e;
	15'h6615: q<=8'h3a;
	15'h6616: q<=8'h00;
	15'h6617: q<=8'h1a;
	15'h6618: q<=8'h16;
	15'h6619: q<=8'h1c;
	15'h661a: q<=8'h16;
	15'h661b: q<=8'h80;
	15'h661c: q<=8'hb8;
	15'h661d: q<=8'h16;
	15'h661e: q<=8'h40;
	15'h661f: q<=8'h32;
	15'h6620: q<=8'h26;
	15'h6621: q<=8'h1c;
	15'h6622: q<=8'h00;
	15'h6623: q<=8'h3a;
	15'h6624: q<=8'h34;
	15'h6625: q<=8'h26;
	15'h6626: q<=8'h2a;
	15'h6627: q<=8'h1e;
	15'h6628: q<=8'hba;
	15'h6629: q<=8'h88;
	15'h662a: q<=8'h16;
	15'h662b: q<=8'h3c;
	15'h662c: q<=8'h3c;
	15'h662d: q<=8'h1e;
	15'h662e: q<=8'h30;
	15'h662f: q<=8'h3c;
	15'h6630: q<=8'h26;
	15'h6631: q<=8'h32;
	15'h6632: q<=8'h30;
	15'h6633: q<=8'h00;
	15'h6634: q<=8'h16;
	15'h6635: q<=8'h3e;
	15'h6636: q<=8'h44;
	15'h6637: q<=8'h00;
	15'h6638: q<=8'h2c;
	15'h6639: q<=8'h16;
	15'h663a: q<=8'h30;
	15'h663b: q<=8'h1a;
	15'h663c: q<=8'h1e;
	15'h663d: q<=8'hba;
	15'h663e: q<=8'h96;
	15'h663f: q<=8'h3a;
	15'h6640: q<=8'h34;
	15'h6641: q<=8'h26;
	15'h6642: q<=8'h3c;
	15'h6643: q<=8'h48;
	15'h6644: q<=8'h1e;
	15'h6645: q<=8'h30;
	15'h6646: q<=8'h00;
	15'h6647: q<=8'h16;
	15'h6648: q<=8'h3e;
	15'h6649: q<=8'h3a;
	15'h664a: q<=8'h42;
	15'h664b: q<=8'h1e;
	15'h664c: q<=8'h26;
	15'h664d: q<=8'h1a;
	15'h664e: q<=8'h24;
	15'h664f: q<=8'h1e;
	15'h6650: q<=8'hb0;
	15'h6651: q<=8'ha0;
	15'h6652: q<=8'h1e;
	15'h6653: q<=8'h40;
	15'h6654: q<=8'h26;
	15'h6655: q<=8'h3c;
	15'h6656: q<=8'h1e;
	15'h6657: q<=8'h00;
	15'h6658: q<=8'h2c;
	15'h6659: q<=8'h16;
	15'h665a: q<=8'h3a;
	15'h665b: q<=8'h00;
	15'h665c: q<=8'h34;
	15'h665d: q<=8'h3e;
	15'h665e: q<=8'h30;
	15'h665f: q<=8'h3c;
	15'h6660: q<=8'h16;
	15'h6661: q<=8'hba;
	15'h6662: q<=8'he0;
	15'h6663: q<=8'h2c;
	15'h6664: q<=8'h1e;
	15'h6665: q<=8'h40;
	15'h6666: q<=8'h1e;
	15'h6667: q<=8'hac;
	15'h6668: q<=8'hda;
	15'h6669: q<=8'h30;
	15'h666a: q<=8'h26;
	15'h666b: q<=8'h40;
	15'h666c: q<=8'h1e;
	15'h666d: q<=8'h16;
	15'h666e: q<=8'hbe;
	15'h666f: q<=8'he2;
	15'h6670: q<=8'h22;
	15'h6671: q<=8'h38;
	15'h6672: q<=8'h16;
	15'h6673: q<=8'h9c;
	15'h6674: q<=8'he0;
	15'h6675: q<=8'h30;
	15'h6676: q<=8'h26;
	15'h6677: q<=8'h40;
	15'h6678: q<=8'h1e;
	15'h6679: q<=8'hac;
	15'h667a: q<=8'hc4;
	15'h667b: q<=8'h3a;
	15'h667c: q<=8'h3e;
	15'h667d: q<=8'h34;
	15'h667e: q<=8'h1e;
	15'h667f: q<=8'h38;
	15'h6680: q<=8'h48;
	15'h6681: q<=8'h16;
	15'h6682: q<=8'h34;
	15'h6683: q<=8'h34;
	15'h6684: q<=8'h1e;
	15'h6685: q<=8'h38;
	15'h6686: q<=8'h00;
	15'h6687: q<=8'h38;
	15'h6688: q<=8'h1e;
	15'h6689: q<=8'h1a;
	15'h668a: q<=8'h24;
	15'h668b: q<=8'h16;
	15'h668c: q<=8'h38;
	15'h668d: q<=8'h22;
	15'h668e: q<=8'h9e;
	15'h668f: q<=8'hcd;
	15'h6690: q<=8'h30;
	15'h6691: q<=8'h1e;
	15'h6692: q<=8'h3e;
	15'h6693: q<=8'h1e;
	15'h6694: q<=8'h38;
	15'h6695: q<=8'h00;
	15'h6696: q<=8'h3a;
	15'h6697: q<=8'h3e;
	15'h6698: q<=8'h34;
	15'h6699: q<=8'h1e;
	15'h669a: q<=8'h38;
	15'h669b: q<=8'h48;
	15'h669c: q<=8'h16;
	15'h669d: q<=8'h34;
	15'h669e: q<=8'h34;
	15'h669f: q<=8'h1e;
	15'h66a0: q<=8'hb8;
	15'h66a1: q<=8'hcd;
	15'h66a2: q<=8'h30;
	15'h66a3: q<=8'h3e;
	15'h66a4: q<=8'h1e;
	15'h66a5: q<=8'h40;
	15'h66a6: q<=8'h32;
	15'h66a7: q<=8'h00;
	15'h66a8: q<=8'h3a;
	15'h66a9: q<=8'h3e;
	15'h66aa: q<=8'h34;
	15'h66ab: q<=8'h1e;
	15'h66ac: q<=8'h38;
	15'h66ad: q<=8'h48;
	15'h66ae: q<=8'h16;
	15'h66af: q<=8'h34;
	15'h66b0: q<=8'h34;
	15'h66b1: q<=8'h1e;
	15'h66b2: q<=8'hb8;
	15'h66b3: q<=8'h31;
	15'h66b4: q<=8'hd0;
	15'h66b5: q<=8'h6d;
	15'h66b6: q<=8'hd0;
	15'h66b7: q<=8'ha9;
	15'h66b8: q<=8'hd0;
	15'h66b9: q<=8'he5;
	15'h66ba: q<=8'hd0;
	15'h66bb: q<=8'had;
	15'h66bc: q<=8'h00;
	15'h66bd: q<=8'h0e;
	15'h66be: q<=8'h85;
	15'h66bf: q<=8'h0a;
	15'h66c0: q<=8'h29;
	15'h66c1: q<=8'h38;
	15'h66c2: q<=8'h4a;
	15'h66c3: q<=8'h4a;
	15'h66c4: q<=8'h4a;
	15'h66c5: q<=8'haa;
	15'h66c6: q<=8'hbd;
	15'h66c7: q<=8'hf7;
	15'h66c8: q<=8'hd6;
	15'h66c9: q<=8'h8d;
	15'h66ca: q<=8'h56;
	15'h66cb: q<=8'h01;
	15'h66cc: q<=8'had;
	15'h66cd: q<=8'h00;
	15'h66ce: q<=8'h0d;
	15'h66cf: q<=8'h49;
	15'h66d0: q<=8'h02;
	15'h66d1: q<=8'h85;
	15'h66d2: q<=8'h09;
	15'h66d3: q<=8'ha5;
	15'h66d4: q<=8'h0a;
	15'h66d5: q<=8'h2a;
	15'h66d6: q<=8'h2a;
	15'h66d7: q<=8'h2a;
	15'h66d8: q<=8'h29;
	15'h66d9: q<=8'h03;
	15'h66da: q<=8'haa;
	15'h66db: q<=8'hbd;
	15'h66dc: q<=8'hff;
	15'h66dd: q<=8'hd6;
	15'h66de: q<=8'h8d;
	15'h66df: q<=8'h58;
	15'h66e0: q<=8'h01;
	15'h66e1: q<=8'ha5;
	15'h66e2: q<=8'h0a;
	15'h66e3: q<=8'h29;
	15'h66e4: q<=8'h06;
	15'h66e5: q<=8'ha8;
	15'h66e6: q<=8'hb9;
	15'h66e7: q<=8'hb3;
	15'h66e8: q<=8'hd6;
	15'h66e9: q<=8'h85;
	15'h66ea: q<=8'hac;
	15'h66eb: q<=8'hb9;
	15'h66ec: q<=8'hb4;
	15'h66ed: q<=8'hd6;
	15'h66ee: q<=8'h85;
	15'h66ef: q<=8'had;
	15'h66f0: q<=8'h20;
	15'h66f1: q<=8'he0;
	15'h66f2: q<=8'hdb;
	15'h66f3: q<=8'h8d;
	15'h66f4: q<=8'h6a;
	15'h66f5: q<=8'h01;
	15'h66f6: q<=8'h60;
	15'h66f7: q<=8'h02;
	15'h66f8: q<=8'h01;
	15'h66f9: q<=8'h03;
	15'h66fa: q<=8'h04;
	15'h66fb: q<=8'h05;
	15'h66fc: q<=8'h06;
	15'h66fd: q<=8'h07;
	15'h66fe: q<=8'h00;
	15'h66ff: q<=8'h03;
	15'h6700: q<=8'h04;
	15'h6701: q<=8'h05;
	15'h6702: q<=8'h02;
	15'h6703: q<=8'h7c;
	15'h6704: q<=8'h48;
	15'h6705: q<=8'h8a;
	15'h6706: q<=8'h48;
	15'h6707: q<=8'h98;
	15'h6708: q<=8'h48;
	15'h6709: q<=8'hd8;
	15'h670a: q<=8'hba;
	15'h670b: q<=8'he0;
	15'h670c: q<=8'hd0;
	15'h670d: q<=8'h90;
	15'h670e: q<=8'h04;
	15'h670f: q<=8'ha5;
	15'h6710: q<=8'h53;
	15'h6711: q<=8'h10;
	15'h6712: q<=8'h04;
	15'h6713: q<=8'h00;
	15'h6714: q<=8'h4c;
	15'h6715: q<=8'h3f;
	15'h6716: q<=8'hd9;
	15'h6717: q<=8'h8d;
	15'h6718: q<=8'h00;
	15'h6719: q<=8'h50;
	15'h671a: q<=8'h8d;
	15'h671b: q<=8'hcb;
	15'h671c: q<=8'h60;
	15'h671d: q<=8'had;
	15'h671e: q<=8'hc8;
	15'h671f: q<=8'h60;
	15'h6720: q<=8'h49;
	15'h6721: q<=8'h0f;
	15'h6722: q<=8'ha8;
	15'h6723: q<=8'h29;
	15'h6724: q<=8'h10;
	15'h6725: q<=8'h8d;
	15'h6726: q<=8'h17;
	15'h6727: q<=8'h01;
	15'h6728: q<=8'h98;
	15'h6729: q<=8'h38;
	15'h672a: q<=8'he5;
	15'h672b: q<=8'h52;
	15'h672c: q<=8'h29;
	15'h672d: q<=8'h0f;
	15'h672e: q<=8'hc9;
	15'h672f: q<=8'h08;
	15'h6730: q<=8'h90;
	15'h6731: q<=8'h02;
	15'h6732: q<=8'h09;
	15'h6733: q<=8'hf0;
	15'h6734: q<=8'h18;
	15'h6735: q<=8'h65;
	15'h6736: q<=8'h50;
	15'h6737: q<=8'h85;
	15'h6738: q<=8'h50;
	15'h6739: q<=8'h84;
	15'h673a: q<=8'h52;
	15'h673b: q<=8'h8d;
	15'h673c: q<=8'hdb;
	15'h673d: q<=8'h60;
	15'h673e: q<=8'hac;
	15'h673f: q<=8'hd8;
	15'h6740: q<=8'h60;
	15'h6741: q<=8'had;
	15'h6742: q<=8'h00;
	15'h6743: q<=8'h0c;
	15'h6744: q<=8'h85;
	15'h6745: q<=8'h08;
	15'h6746: q<=8'ha5;
	15'h6747: q<=8'h4c;
	15'h6748: q<=8'h84;
	15'h6749: q<=8'h4c;
	15'h674a: q<=8'ha8;
	15'h674b: q<=8'h25;
	15'h674c: q<=8'h4c;
	15'h674d: q<=8'h05;
	15'h674e: q<=8'h4d;
	15'h674f: q<=8'h85;
	15'h6750: q<=8'h4d;
	15'h6751: q<=8'h98;
	15'h6752: q<=8'h05;
	15'h6753: q<=8'h4c;
	15'h6754: q<=8'h25;
	15'h6755: q<=8'h4d;
	15'h6756: q<=8'h85;
	15'h6757: q<=8'h4d;
	15'h6758: q<=8'ha8;
	15'h6759: q<=8'h45;
	15'h675a: q<=8'h4f;
	15'h675b: q<=8'h25;
	15'h675c: q<=8'h4d;
	15'h675d: q<=8'h05;
	15'h675e: q<=8'h4e;
	15'h675f: q<=8'h85;
	15'h6760: q<=8'h4e;
	15'h6761: q<=8'h84;
	15'h6762: q<=8'h4f;
	15'h6763: q<=8'ha5;
	15'h6764: q<=8'hb4;
	15'h6765: q<=8'ha4;
	15'h6766: q<=8'h13;
	15'h6767: q<=8'h10;
	15'h6768: q<=8'h02;
	15'h6769: q<=8'h09;
	15'h676a: q<=8'h04;
	15'h676b: q<=8'ha4;
	15'h676c: q<=8'h14;
	15'h676d: q<=8'h10;
	15'h676e: q<=8'h02;
	15'h676f: q<=8'h09;
	15'h6770: q<=8'h02;
	15'h6771: q<=8'ha4;
	15'h6772: q<=8'h15;
	15'h6773: q<=8'h10;
	15'h6774: q<=8'h02;
	15'h6775: q<=8'h09;
	15'h6776: q<=8'h01;
	15'h6777: q<=8'h8d;
	15'h6778: q<=8'h00;
	15'h6779: q<=8'h40;
	15'h677a: q<=8'ha6;
	15'h677b: q<=8'h3e;
	15'h677c: q<=8'he8;
	15'h677d: q<=8'ha4;
	15'h677e: q<=8'h05;
	15'h677f: q<=8'hd0;
	15'h6780: q<=8'h10;
	15'h6781: q<=8'ha2;
	15'h6782: q<=8'h00;
	15'h6783: q<=8'ha4;
	15'h6784: q<=8'h07;
	15'h6785: q<=8'hc0;
	15'h6786: q<=8'h40;
	15'h6787: q<=8'h90;
	15'h6788: q<=8'h08;
	15'h6789: q<=8'ha6;
	15'h678a: q<=8'h06;
	15'h678b: q<=8'he0;
	15'h678c: q<=8'h02;
	15'h678d: q<=8'h90;
	15'h678e: q<=8'h02;
	15'h678f: q<=8'ha2;
	15'h6790: q<=8'h03;
	15'h6791: q<=8'hbd;
	15'h6792: q<=8'hdd;
	15'h6793: q<=8'hd7;
	15'h6794: q<=8'h45;
	15'h6795: q<=8'ha1;
	15'h6796: q<=8'h29;
	15'h6797: q<=8'h03;
	15'h6798: q<=8'h45;
	15'h6799: q<=8'ha1;
	15'h679a: q<=8'h85;
	15'h679b: q<=8'ha1;
	15'h679c: q<=8'h8d;
	15'h679d: q<=8'he0;
	15'h679e: q<=8'h60;
	15'h679f: q<=8'h20;
	15'h67a0: q<=8'h24;
	15'h67a1: q<=8'hcf;
	15'h67a2: q<=8'h20;
	15'h67a3: q<=8'h0a;
	15'h67a4: q<=8'hcd;
	15'h67a5: q<=8'he6;
	15'h67a6: q<=8'h53;
	15'h67a7: q<=8'he6;
	15'h67a8: q<=8'h07;
	15'h67a9: q<=8'hd0;
	15'h67aa: q<=8'h1e;
	15'h67ab: q<=8'hee;
	15'h67ac: q<=8'h06;
	15'h67ad: q<=8'h04;
	15'h67ae: q<=8'hd0;
	15'h67af: q<=8'h08;
	15'h67b0: q<=8'hee;
	15'h67b1: q<=8'h07;
	15'h67b2: q<=8'h04;
	15'h67b3: q<=8'hd0;
	15'h67b4: q<=8'h03;
	15'h67b5: q<=8'hee;
	15'h67b6: q<=8'h08;
	15'h67b7: q<=8'h04;
	15'h67b8: q<=8'h24;
	15'h67b9: q<=8'h05;
	15'h67ba: q<=8'h50;
	15'h67bb: q<=8'h0d;
	15'h67bc: q<=8'hee;
	15'h67bd: q<=8'h09;
	15'h67be: q<=8'h04;
	15'h67bf: q<=8'hd0;
	15'h67c0: q<=8'h08;
	15'h67c1: q<=8'hee;
	15'h67c2: q<=8'h0a;
	15'h67c3: q<=8'h04;
	15'h67c4: q<=8'hd0;
	15'h67c5: q<=8'h03;
	15'h67c6: q<=8'hee;
	15'h67c7: q<=8'h0b;
	15'h67c8: q<=8'h04;
	15'h67c9: q<=8'h2c;
	15'h67ca: q<=8'h00;
	15'h67cb: q<=8'h0c;
	15'h67cc: q<=8'h50;
	15'h67cd: q<=8'h09;
	15'h67ce: q<=8'hee;
	15'h67cf: q<=8'h33;
	15'h67d0: q<=8'h01;
	15'h67d1: q<=8'h8d;
	15'h67d2: q<=8'h00;
	15'h67d3: q<=8'h58;
	15'h67d4: q<=8'h8d;
	15'h67d5: q<=8'h00;
	15'h67d6: q<=8'h48;
	15'h67d7: q<=8'h68;
	15'h67d8: q<=8'ha8;
	15'h67d9: q<=8'h68;
	15'h67da: q<=8'haa;
	15'h67db: q<=8'h68;
	15'h67dc: q<=8'h40;
	15'h67dd: q<=8'hff;
	15'h67de: q<=8'hfd;
	15'h67df: q<=8'hfe;
	15'h67e0: q<=8'hfc;
	15'h67e1: q<=8'ha9;
	15'h67e2: q<=8'h00;
	15'h67e3: q<=8'h85;
	15'h67e4: q<=8'h05;
	15'h67e5: q<=8'ha9;
	15'h67e6: q<=8'h02;
	15'h67e7: q<=8'h85;
	15'h67e8: q<=8'h01;
	15'h67e9: q<=8'had;
	15'h67ea: q<=8'hca;
	15'h67eb: q<=8'h01;
	15'h67ec: q<=8'hd0;
	15'h67ed: q<=8'h15;
	15'h67ee: q<=8'had;
	15'h67ef: q<=8'h00;
	15'h67f0: q<=8'h0c;
	15'h67f1: q<=8'h29;
	15'h67f2: q<=8'h10;
	15'h67f3: q<=8'hf0;
	15'h67f4: q<=8'h0e;
	15'h67f5: q<=8'ha9;
	15'h67f6: q<=8'h00;
	15'h67f7: q<=8'h85;
	15'h67f8: q<=8'h00;
	15'h67f9: q<=8'had;
	15'h67fa: q<=8'hc9;
	15'h67fb: q<=8'h01;
	15'h67fc: q<=8'h29;
	15'h67fd: q<=8'h03;
	15'h67fe: q<=8'hf0;
	15'h67ff: q<=8'h03;
	15'h6800: q<=8'h20;
	15'h6801: q<=8'hac;
	15'h6802: q<=8'hab;
	15'h6803: q<=8'h60;
	15'h6804: q<=8'h20;
	15'h6805: q<=8'hbb;
	15'h6806: q<=8'hd6;
	15'h6807: q<=8'h20;
	15'h6808: q<=8'ha8;
	15'h6809: q<=8'haa;
	15'h680a: q<=8'h20;
	15'h680b: q<=8'h0d;
	15'h680c: q<=8'hdd;
	15'h680d: q<=8'h20;
	15'h680e: q<=8'h41;
	15'h680f: q<=8'hdd;
	15'h6810: q<=8'had;
	15'h6811: q<=8'h58;
	15'h6812: q<=8'h01;
	15'h6813: q<=8'h85;
	15'h6814: q<=8'h37;
	15'h6815: q<=8'h20;
	15'h6816: q<=8'h53;
	15'h6817: q<=8'hdf;
	15'h6818: q<=8'ha9;
	15'h6819: q<=8'he8;
	15'h681a: q<=8'ha2;
	15'h681b: q<=8'hc0;
	15'h681c: q<=8'h20;
	15'h681d: q<=8'h75;
	15'h681e: q<=8'hdf;
	15'h681f: q<=8'ha9;
	15'h6820: q<=8'h32;
	15'h6821: q<=8'ha2;
	15'h6822: q<=8'h6c;
	15'h6823: q<=8'h20;
	15'h6824: q<=8'h39;
	15'h6825: q<=8'hdf;
	15'h6826: q<=8'hc6;
	15'h6827: q<=8'h37;
	15'h6828: q<=8'hd0;
	15'h6829: q<=8'hf5;
	15'h682a: q<=8'had;
	15'h682b: q<=8'h6a;
	15'h682c: q<=8'h01;
	15'h682d: q<=8'h29;
	15'h682e: q<=8'h03;
	15'h682f: q<=8'h0a;
	15'h6830: q<=8'ha8;
	15'h6831: q<=8'hb9;
	15'h6832: q<=8'h1f;
	15'h6833: q<=8'h3f;
	15'h6834: q<=8'hbe;
	15'h6835: q<=8'h1e;
	15'h6836: q<=8'h3f;
	15'h6837: q<=8'h20;
	15'h6838: q<=8'h39;
	15'h6839: q<=8'hdf;
	15'h683a: q<=8'had;
	15'h683b: q<=8'h00;
	15'h683c: q<=8'h02;
	15'h683d: q<=8'h20;
	15'h683e: q<=8'hce;
	15'h683f: q<=8'had;
	15'h6840: q<=8'h8d;
	15'h6841: q<=8'h00;
	15'h6842: q<=8'h02;
	15'h6843: q<=8'h29;
	15'h6844: q<=8'h06;
	15'h6845: q<=8'h48;
	15'h6846: q<=8'ha8;
	15'h6847: q<=8'hb9;
	15'h6848: q<=8'h17;
	15'h6849: q<=8'h3f;
	15'h684a: q<=8'hbe;
	15'h684b: q<=8'h16;
	15'h684c: q<=8'h3f;
	15'h684d: q<=8'h20;
	15'h684e: q<=8'h39;
	15'h684f: q<=8'hdf;
	15'h6850: q<=8'h68;
	15'h6851: q<=8'h4a;
	15'h6852: q<=8'haa;
	15'h6853: q<=8'ha5;
	15'h6854: q<=8'h4d;
	15'h6855: q<=8'h3d;
	15'h6856: q<=8'hb6;
	15'h6857: q<=8'hd8;
	15'h6858: q<=8'hdd;
	15'h6859: q<=8'hb6;
	15'h685a: q<=8'hd8;
	15'h685b: q<=8'hd0;
	15'h685c: q<=8'h1a;
	15'h685d: q<=8'hca;
	15'h685e: q<=8'hca;
	15'h685f: q<=8'h10;
	15'h6860: q<=8'h03;
	15'h6861: q<=8'h4c;
	15'h6862: q<=8'h3f;
	15'h6863: q<=8'hd9;
	15'h6864: q<=8'hd0;
	15'h6865: q<=8'h06;
	15'h6866: q<=8'h20;
	15'h6867: q<=8'he9;
	15'h6868: q<=8'hdd;
	15'h6869: q<=8'hb8;
	15'h686a: q<=8'h50;
	15'h686b: q<=8'h0b;
	15'h686c: q<=8'h20;
	15'h686d: q<=8'hed;
	15'h686e: q<=8'hdd;
	15'h686f: q<=8'had;
	15'h6870: q<=8'hc9;
	15'h6871: q<=8'h01;
	15'h6872: q<=8'h09;
	15'h6873: q<=8'h03;
	15'h6874: q<=8'h8d;
	15'h6875: q<=8'hc9;
	15'h6876: q<=8'h01;
	15'h6877: q<=8'had;
	15'h6878: q<=8'hca;
	15'h6879: q<=8'h01;
	15'h687a: q<=8'h2d;
	15'h687b: q<=8'hc6;
	15'h687c: q<=8'h01;
	15'h687d: q<=8'hf0;
	15'h687e: q<=8'h07;
	15'h687f: q<=8'ha9;
	15'h6880: q<=8'h34;
	15'h6881: q<=8'ha2;
	15'h6882: q<=8'h6e;
	15'h6883: q<=8'h20;
	15'h6884: q<=8'h39;
	15'h6885: q<=8'hdf;
	15'h6886: q<=8'h20;
	15'h6887: q<=8'h53;
	15'h6888: q<=8'hdf;
	15'h6889: q<=8'ha5;
	15'h688a: q<=8'h09;
	15'h688b: q<=8'h29;
	15'h688c: q<=8'h1c;
	15'h688d: q<=8'h4a;
	15'h688e: q<=8'h4a;
	15'h688f: q<=8'haa;
	15'h6890: q<=8'hbd;
	15'h6891: q<=8'hba;
	15'h6892: q<=8'hd8;
	15'h6893: q<=8'ha0;
	15'h6894: q<=8'hee;
	15'h6895: q<=8'ha2;
	15'h6896: q<=8'h1b;
	15'h6897: q<=8'h20;
	15'h6898: q<=8'ha9;
	15'h6899: q<=8'hd8;
	15'h689a: q<=8'ha5;
	15'h689b: q<=8'h09;
	15'h689c: q<=8'h4a;
	15'h689d: q<=8'h4a;
	15'h689e: q<=8'h4a;
	15'h689f: q<=8'h4a;
	15'h68a0: q<=8'h4a;
	15'h68a1: q<=8'haa;
	15'h68a2: q<=8'hbd;
	15'h68a3: q<=8'hc2;
	15'h68a4: q<=8'hd8;
	15'h68a5: q<=8'ha0;
	15'h68a6: q<=8'h32;
	15'h68a7: q<=8'ha2;
	15'h68a8: q<=8'hf8;
	15'h68a9: q<=8'h85;
	15'h68aa: q<=8'h29;
	15'h68ab: q<=8'h98;
	15'h68ac: q<=8'h20;
	15'h68ad: q<=8'h75;
	15'h68ae: q<=8'hdf;
	15'h68af: q<=8'ha9;
	15'h68b0: q<=8'h29;
	15'h68b1: q<=8'ha0;
	15'h68b2: q<=8'h01;
	15'h68b3: q<=8'h4c;
	15'h68b4: q<=8'hb1;
	15'h68b5: q<=8'hdf;
	15'h68b6: q<=8'h18;
	15'h68b7: q<=8'h18;
	15'h68b8: q<=8'h30;
	15'h68b9: q<=8'h50;
	15'h68ba: q<=8'h11;
	15'h68bb: q<=8'h14;
	15'h68bc: q<=8'h15;
	15'h68bd: q<=8'h16;
	15'h68be: q<=8'h21;
	15'h68bf: q<=8'h24;
	15'h68c0: q<=8'h25;
	15'h68c1: q<=8'h26;
	15'h68c2: q<=8'h00;
	15'h68c3: q<=8'h12;
	15'h68c4: q<=8'h14;
	15'h68c5: q<=8'h24;
	15'h68c6: q<=8'h15;
	15'h68c7: q<=8'h13;
	15'h68c8: q<=8'h00;
	15'h68c9: q<=8'h00;
	15'h68ca: q<=8'ha8;
	15'h68cb: q<=8'ha9;
	15'h68cc: q<=8'h00;
	15'h68cd: q<=8'h84;
	15'h68ce: q<=8'h79;
	15'h68cf: q<=8'h4a;
	15'h68d0: q<=8'h4a;
	15'h68d1: q<=8'h0a;
	15'h68d2: q<=8'haa;
	15'h68d3: q<=8'h98;
	15'h68d4: q<=8'h29;
	15'h68d5: q<=8'h0f;
	15'h68d6: q<=8'hd0;
	15'h68d7: q<=8'h01;
	15'h68d8: q<=8'he8;
	15'h68d9: q<=8'h9a;
	15'h68da: q<=8'ha9;
	15'h68db: q<=8'ha2;
	15'h68dc: q<=8'h8d;
	15'h68dd: q<=8'hc1;
	15'h68de: q<=8'h60;
	15'h68df: q<=8'hba;
	15'h68e0: q<=8'hd0;
	15'h68e1: q<=8'h07;
	15'h68e2: q<=8'ha9;
	15'h68e3: q<=8'h60;
	15'h68e4: q<=8'ha0;
	15'h68e5: q<=8'h09;
	15'h68e6: q<=8'hb8;
	15'h68e7: q<=8'h50;
	15'h68e8: q<=8'h04;
	15'h68e9: q<=8'ha9;
	15'h68ea: q<=8'hc0;
	15'h68eb: q<=8'ha0;
	15'h68ec: q<=8'h01;
	15'h68ed: q<=8'h8d;
	15'h68ee: q<=8'hc0;
	15'h68ef: q<=8'h60;
	15'h68f0: q<=8'ha9;
	15'h68f1: q<=8'h03;
	15'h68f2: q<=8'h8d;
	15'h68f3: q<=8'he0;
	15'h68f4: q<=8'h60;
	15'h68f5: q<=8'ha2;
	15'h68f6: q<=8'h00;
	15'h68f7: q<=8'h2c;
	15'h68f8: q<=8'h00;
	15'h68f9: q<=8'h0c;
	15'h68fa: q<=8'h30;
	15'h68fb: q<=8'hfb;
	15'h68fc: q<=8'h2c;
	15'h68fd: q<=8'h00;
	15'h68fe: q<=8'h0c;
	15'h68ff: q<=8'h10;
	15'h6900: q<=8'hfb;
	15'h6901: q<=8'h8d;
	15'h6902: q<=8'h00;
	15'h6903: q<=8'h50;
	15'h6904: q<=8'hca;
	15'h6905: q<=8'hd0;
	15'h6906: q<=8'hf0;
	15'h6907: q<=8'h88;
	15'h6908: q<=8'hd0;
	15'h6909: q<=8'hed;
	15'h690a: q<=8'h8e;
	15'h690b: q<=8'hc1;
	15'h690c: q<=8'h60;
	15'h690d: q<=8'ha9;
	15'h690e: q<=8'h00;
	15'h690f: q<=8'h8d;
	15'h6910: q<=8'he0;
	15'h6911: q<=8'h60;
	15'h6912: q<=8'ha0;
	15'h6913: q<=8'h09;
	15'h6914: q<=8'h2c;
	15'h6915: q<=8'h00;
	15'h6916: q<=8'h0c;
	15'h6917: q<=8'h30;
	15'h6918: q<=8'hfb;
	15'h6919: q<=8'h2c;
	15'h691a: q<=8'h00;
	15'h691b: q<=8'h0c;
	15'h691c: q<=8'h10;
	15'h691d: q<=8'hfb;
	15'h691e: q<=8'h8d;
	15'h691f: q<=8'h00;
	15'h6920: q<=8'h50;
	15'h6921: q<=8'hca;
	15'h6922: q<=8'hd0;
	15'h6923: q<=8'hf0;
	15'h6924: q<=8'h88;
	15'h6925: q<=8'hd0;
	15'h6926: q<=8'hed;
	15'h6927: q<=8'hba;
	15'h6928: q<=8'hca;
	15'h6929: q<=8'h9a;
	15'h692a: q<=8'h10;
	15'h692b: q<=8'hae;
	15'h692c: q<=8'h4c;
	15'h692d: q<=8'h0a;
	15'h692e: q<=8'hda;
	15'h692f: q<=8'h51;
	15'h6930: q<=8'h00;
	15'h6931: q<=8'ha8;
	15'h6932: q<=8'ha5;
	15'h6933: q<=8'h01;
	15'h6934: q<=8'hc9;
	15'h6935: q<=8'h20;
	15'h6936: q<=8'h90;
	15'h6937: q<=8'h02;
	15'h6938: q<=8'he9;
	15'h6939: q<=8'h18;
	15'h693a: q<=8'h29;
	15'h693b: q<=8'h1f;
	15'h693c: q<=8'h4c;
	15'h693d: q<=8'hcd;
	15'h693e: q<=8'hd8;
	15'h693f: q<=8'h78;
	15'h6940: q<=8'h8d;
	15'h6941: q<=8'h00;
	15'h6942: q<=8'h50;
	15'h6943: q<=8'h8d;
	15'h6944: q<=8'h00;
	15'h6945: q<=8'h58;
	15'h6946: q<=8'ha2;
	15'h6947: q<=8'hff;
	15'h6948: q<=8'h9a;
	15'h6949: q<=8'hd8;
	15'h694a: q<=8'he8;
	15'h694b: q<=8'h8a;
	15'h694c: q<=8'ha8;
	15'h694d: q<=8'h84;
	15'h694e: q<=8'h00;
	15'h694f: q<=8'h86;
	15'h6950: q<=8'h01;
	15'h6951: q<=8'ha0;
	15'h6952: q<=8'h00;
	15'h6953: q<=8'h91;
	15'h6954: q<=8'h00;
	15'h6955: q<=8'hc8;
	15'h6956: q<=8'hd0;
	15'h6957: q<=8'hfb;
	15'h6958: q<=8'he8;
	15'h6959: q<=8'he0;
	15'h695a: q<=8'h08;
	15'h695b: q<=8'hd0;
	15'h695c: q<=8'h02;
	15'h695d: q<=8'ha2;
	15'h695e: q<=8'h20;
	15'h695f: q<=8'he0;
	15'h6960: q<=8'h30;
	15'h6961: q<=8'h8d;
	15'h6962: q<=8'h00;
	15'h6963: q<=8'h50;
	15'h6964: q<=8'h90;
	15'h6965: q<=8'he7;
	15'h6966: q<=8'h85;
	15'h6967: q<=8'h01;
	15'h6968: q<=8'h8d;
	15'h6969: q<=8'he0;
	15'h696a: q<=8'h60;
	15'h696b: q<=8'h8d;
	15'h696c: q<=8'hcf;
	15'h696d: q<=8'h60;
	15'h696e: q<=8'h8d;
	15'h696f: q<=8'hdf;
	15'h6970: q<=8'h60;
	15'h6971: q<=8'ha2;
	15'h6972: q<=8'h07;
	15'h6973: q<=8'h8e;
	15'h6974: q<=8'hcf;
	15'h6975: q<=8'h60;
	15'h6976: q<=8'h8e;
	15'h6977: q<=8'hdf;
	15'h6978: q<=8'h60;
	15'h6979: q<=8'he8;
	15'h697a: q<=8'h9d;
	15'h697b: q<=8'hc0;
	15'h697c: q<=8'h60;
	15'h697d: q<=8'h9d;
	15'h697e: q<=8'hd0;
	15'h697f: q<=8'h60;
	15'h6980: q<=8'hca;
	15'h6981: q<=8'h10;
	15'h6982: q<=8'hf7;
	15'h6983: q<=8'had;
	15'h6984: q<=8'h00;
	15'h6985: q<=8'h0c;
	15'h6986: q<=8'h29;
	15'h6987: q<=8'h10;
	15'h6988: q<=8'hf0;
	15'h6989: q<=8'h1f;
	15'h698a: q<=8'h8d;
	15'h698b: q<=8'h00;
	15'h698c: q<=8'h50;
	15'h698d: q<=8'hce;
	15'h698e: q<=8'h00;
	15'h698f: q<=8'h01;
	15'h6990: q<=8'hd0;
	15'h6991: q<=8'hf8;
	15'h6992: q<=8'hce;
	15'h6993: q<=8'h01;
	15'h6994: q<=8'h01;
	15'h6995: q<=8'hd0;
	15'h6996: q<=8'hf3;
	15'h6997: q<=8'ha9;
	15'h6998: q<=8'h10;
	15'h6999: q<=8'h85;
	15'h699a: q<=8'hb4;
	15'h699b: q<=8'h20;
	15'h699c: q<=8'h11;
	15'h699d: q<=8'hde;
	15'h699e: q<=8'h20;
	15'h699f: q<=8'hac;
	15'h69a0: q<=8'hab;
	15'h69a1: q<=8'h20;
	15'h69a2: q<=8'h6e;
	15'h69a3: q<=8'hc1;
	15'h69a4: q<=8'h58;
	15'h69a5: q<=8'h4c;
	15'h69a6: q<=8'ha0;
	15'h69a7: q<=8'hc7;
	15'h69a8: q<=8'ha0;
	15'h69a9: q<=8'ha2;
	15'h69aa: q<=8'h11;
	15'h69ab: q<=8'h9a;
	15'h69ac: q<=8'ha0;
	15'h69ad: q<=8'h00;
	15'h69ae: q<=8'hba;
	15'h69af: q<=8'h96;
	15'h69b0: q<=8'h00;
	15'h69b1: q<=8'ha2;
	15'h69b2: q<=8'h01;
	15'h69b3: q<=8'hc8;
	15'h69b4: q<=8'hb9;
	15'h69b5: q<=8'h00;
	15'h69b6: q<=8'h00;
	15'h69b7: q<=8'hf0;
	15'h69b8: q<=8'h03;
	15'h69b9: q<=8'h4c;
	15'h69ba: q<=8'hca;
	15'h69bb: q<=8'hd8;
	15'h69bc: q<=8'he8;
	15'h69bd: q<=8'hd0;
	15'h69be: q<=8'hf4;
	15'h69bf: q<=8'hba;
	15'h69c0: q<=8'h8a;
	15'h69c1: q<=8'h8d;
	15'h69c2: q<=8'h00;
	15'h69c3: q<=8'h50;
	15'h69c4: q<=8'hc8;
	15'h69c5: q<=8'h59;
	15'h69c6: q<=8'h00;
	15'h69c7: q<=8'h00;
	15'h69c8: q<=8'hd0;
	15'h69c9: q<=8'hef;
	15'h69ca: q<=8'h99;
	15'h69cb: q<=8'h00;
	15'h69cc: q<=8'h00;
	15'h69cd: q<=8'hc8;
	15'h69ce: q<=8'hd0;
	15'h69cf: q<=8'hde;
	15'h69d0: q<=8'hba;
	15'h69d1: q<=8'h8a;
	15'h69d2: q<=8'h0a;
	15'h69d3: q<=8'haa;
	15'h69d4: q<=8'h90;
	15'h69d5: q<=8'hd5;
	15'h69d6: q<=8'ha0;
	15'h69d7: q<=8'h00;
	15'h69d8: q<=8'ha2;
	15'h69d9: q<=8'h01;
	15'h69da: q<=8'h84;
	15'h69db: q<=8'h00;
	15'h69dc: q<=8'h86;
	15'h69dd: q<=8'h01;
	15'h69de: q<=8'ha0;
	15'h69df: q<=8'h00;
	15'h69e0: q<=8'hb1;
	15'h69e1: q<=8'h00;
	15'h69e2: q<=8'hf0;
	15'h69e3: q<=8'h03;
	15'h69e4: q<=8'h4c;
	15'h69e5: q<=8'h31;
	15'h69e6: q<=8'hd9;
	15'h69e7: q<=8'ha9;
	15'h69e8: q<=8'h11;
	15'h69e9: q<=8'h91;
	15'h69ea: q<=8'h00;
	15'h69eb: q<=8'hd1;
	15'h69ec: q<=8'h00;
	15'h69ed: q<=8'hf0;
	15'h69ee: q<=8'h03;
	15'h69ef: q<=8'h4c;
	15'h69f0: q<=8'h2f;
	15'h69f1: q<=8'hd9;
	15'h69f2: q<=8'h0a;
	15'h69f3: q<=8'h90;
	15'h69f4: q<=8'hf4;
	15'h69f5: q<=8'ha9;
	15'h69f6: q<=8'h00;
	15'h69f7: q<=8'h91;
	15'h69f8: q<=8'h00;
	15'h69f9: q<=8'hc8;
	15'h69fa: q<=8'hd0;
	15'h69fb: q<=8'he4;
	15'h69fc: q<=8'h8d;
	15'h69fd: q<=8'h00;
	15'h69fe: q<=8'h50;
	15'h69ff: q<=8'he8;
	15'h6a00: q<=8'he0;
	15'h6a01: q<=8'h08;
	15'h6a02: q<=8'hd0;
	15'h6a03: q<=8'h02;
	15'h6a04: q<=8'ha2;
	15'h6a05: q<=8'h20;
	15'h6a06: q<=8'he0;
	15'h6a07: q<=8'h30;
	15'h6a08: q<=8'h90;
	15'h6a09: q<=8'hd0;
	15'h6a0a: q<=8'ha9;
	15'h6a0b: q<=8'h00;
	15'h6a0c: q<=8'ha8;
	15'h6a0d: q<=8'haa;
	15'h6a0e: q<=8'h85;
	15'h6a0f: q<=8'h3b;
	15'h6a10: q<=8'ha9;
	15'h6a11: q<=8'h30;
	15'h6a12: q<=8'h85;
	15'h6a13: q<=8'h3c;
	15'h6a14: q<=8'ha9;
	15'h6a15: q<=8'h08;
	15'h6a16: q<=8'h85;
	15'h6a17: q<=8'h38;
	15'h6a18: q<=8'h8a;
	15'h6a19: q<=8'h51;
	15'h6a1a: q<=8'h3b;
	15'h6a1b: q<=8'hc8;
	15'h6a1c: q<=8'hd0;
	15'h6a1d: q<=8'hfb;
	15'h6a1e: q<=8'he6;
	15'h6a1f: q<=8'h3c;
	15'h6a20: q<=8'h8d;
	15'h6a21: q<=8'h00;
	15'h6a22: q<=8'h50;
	15'h6a23: q<=8'hc6;
	15'h6a24: q<=8'h38;
	15'h6a25: q<=8'hd0;
	15'h6a26: q<=8'hf2;
	15'h6a27: q<=8'h95;
	15'h6a28: q<=8'h7d;
	15'h6a29: q<=8'he8;
	15'h6a2a: q<=8'he0;
	15'h6a2b: q<=8'h02;
	15'h6a2c: q<=8'hd0;
	15'h6a2d: q<=8'h04;
	15'h6a2e: q<=8'ha9;
	15'h6a2f: q<=8'h90;
	15'h6a30: q<=8'h85;
	15'h6a31: q<=8'h3c;
	15'h6a32: q<=8'he0;
	15'h6a33: q<=8'h0c;
	15'h6a34: q<=8'h90;
	15'h6a35: q<=8'hde;
	15'h6a36: q<=8'ha5;
	15'h6a37: q<=8'h7d;
	15'h6a38: q<=8'hf0;
	15'h6a39: q<=8'h0a;
	15'h6a3a: q<=8'ha9;
	15'h6a3b: q<=8'h40;
	15'h6a3c: q<=8'ha2;
	15'h6a3d: q<=8'ha4;
	15'h6a3e: q<=8'h8d;
	15'h6a3f: q<=8'hc4;
	15'h6a40: q<=8'h60;
	15'h6a41: q<=8'h8e;
	15'h6a42: q<=8'hc5;
	15'h6a43: q<=8'h60;
	15'h6a44: q<=8'ha2;
	15'h6a45: q<=8'h05;
	15'h6a46: q<=8'had;
	15'h6a47: q<=8'hca;
	15'h6a48: q<=8'h60;
	15'h6a49: q<=8'hcd;
	15'h6a4a: q<=8'hca;
	15'h6a4b: q<=8'h60;
	15'h6a4c: q<=8'hd0;
	15'h6a4d: q<=8'h05;
	15'h6a4e: q<=8'hca;
	15'h6a4f: q<=8'h10;
	15'h6a50: q<=8'hf8;
	15'h6a51: q<=8'h85;
	15'h6a52: q<=8'h7a;
	15'h6a53: q<=8'ha2;
	15'h6a54: q<=8'h05;
	15'h6a55: q<=8'had;
	15'h6a56: q<=8'hda;
	15'h6a57: q<=8'h60;
	15'h6a58: q<=8'hcd;
	15'h6a59: q<=8'hda;
	15'h6a5a: q<=8'h60;
	15'h6a5b: q<=8'hd0;
	15'h6a5c: q<=8'h05;
	15'h6a5d: q<=8'hca;
	15'h6a5e: q<=8'h10;
	15'h6a5f: q<=8'hf8;
	15'h6a60: q<=8'h85;
	15'h6a61: q<=8'h7b;
	15'h6a62: q<=8'h20;
	15'h6a63: q<=8'h11;
	15'h6a64: q<=8'hde;
	15'h6a65: q<=8'ha0;
	15'h6a66: q<=8'h02;
	15'h6a67: q<=8'had;
	15'h6a68: q<=8'hc9;
	15'h6a69: q<=8'h01;
	15'h6a6a: q<=8'hf0;
	15'h6a6b: q<=8'h0a;
	15'h6a6c: q<=8'h85;
	15'h6a6d: q<=8'h7c;
	15'h6a6e: q<=8'h20;
	15'h6a6f: q<=8'hf1;
	15'h6a70: q<=8'hdd;
	15'h6a71: q<=8'ha0;
	15'h6a72: q<=8'h00;
	15'h6a73: q<=8'h8c;
	15'h6a74: q<=8'hc9;
	15'h6a75: q<=8'h01;
	15'h6a76: q<=8'h84;
	15'h6a77: q<=8'h00;
	15'h6a78: q<=8'ha2;
	15'h6a79: q<=8'h07;
	15'h6a7a: q<=8'hbd;
	15'h6a7b: q<=8'hf9;
	15'h6a7c: q<=8'hda;
	15'h6a7d: q<=8'h9d;
	15'h6a7e: q<=8'h00;
	15'h6a7f: q<=8'h08;
	15'h6a80: q<=8'hca;
	15'h6a81: q<=8'h10;
	15'h6a82: q<=8'hf7;
	15'h6a83: q<=8'ha9;
	15'h6a84: q<=8'h00;
	15'h6a85: q<=8'h8d;
	15'h6a86: q<=8'he0;
	15'h6a87: q<=8'h60;
	15'h6a88: q<=8'ha9;
	15'h6a89: q<=8'h10;
	15'h6a8a: q<=8'h8d;
	15'h6a8b: q<=8'h00;
	15'h6a8c: q<=8'h40;
	15'h6a8d: q<=8'ha0;
	15'h6a8e: q<=8'h04;
	15'h6a8f: q<=8'ha2;
	15'h6a90: q<=8'h14;
	15'h6a91: q<=8'h2c;
	15'h6a92: q<=8'h00;
	15'h6a93: q<=8'h0c;
	15'h6a94: q<=8'h10;
	15'h6a95: q<=8'hfb;
	15'h6a96: q<=8'h2c;
	15'h6a97: q<=8'h00;
	15'h6a98: q<=8'h0c;
	15'h6a99: q<=8'h30;
	15'h6a9a: q<=8'hfb;
	15'h6a9b: q<=8'hca;
	15'h6a9c: q<=8'h10;
	15'h6a9d: q<=8'hf3;
	15'h6a9e: q<=8'h88;
	15'h6a9f: q<=8'h30;
	15'h6aa0: q<=8'h08;
	15'h6aa1: q<=8'h8d;
	15'h6aa2: q<=8'h00;
	15'h6aa3: q<=8'h50;
	15'h6aa4: q<=8'h2c;
	15'h6aa5: q<=8'h00;
	15'h6aa6: q<=8'h0c;
	15'h6aa7: q<=8'h50;
	15'h6aa8: q<=8'he6;
	15'h6aa9: q<=8'h8d;
	15'h6aaa: q<=8'h00;
	15'h6aab: q<=8'h58;
	15'h6aac: q<=8'ha9;
	15'h6aad: q<=8'h00;
	15'h6aae: q<=8'h85;
	15'h6aaf: q<=8'h74;
	15'h6ab0: q<=8'ha9;
	15'h6ab1: q<=8'h20;
	15'h6ab2: q<=8'h85;
	15'h6ab3: q<=8'h75;
	15'h6ab4: q<=8'h8d;
	15'h6ab5: q<=8'hcb;
	15'h6ab6: q<=8'h60;
	15'h6ab7: q<=8'had;
	15'h6ab8: q<=8'hc8;
	15'h6ab9: q<=8'h60;
	15'h6aba: q<=8'h85;
	15'h6abb: q<=8'h52;
	15'h6abc: q<=8'h29;
	15'h6abd: q<=8'h0f;
	15'h6abe: q<=8'h85;
	15'h6abf: q<=8'h50;
	15'h6ac0: q<=8'had;
	15'h6ac1: q<=8'h00;
	15'h6ac2: q<=8'h0c;
	15'h6ac3: q<=8'h49;
	15'h6ac4: q<=8'hff;
	15'h6ac5: q<=8'h29;
	15'h6ac6: q<=8'h2f;
	15'h6ac7: q<=8'h85;
	15'h6ac8: q<=8'h4e;
	15'h6ac9: q<=8'h29;
	15'h6aca: q<=8'h28;
	15'h6acb: q<=8'hf0;
	15'h6acc: q<=8'h0b;
	15'h6acd: q<=8'h06;
	15'h6ace: q<=8'h4c;
	15'h6acf: q<=8'h90;
	15'h6ad0: q<=8'h04;
	15'h6ad1: q<=8'he6;
	15'h6ad2: q<=8'h00;
	15'h6ad3: q<=8'he6;
	15'h6ad4: q<=8'h00;
	15'h6ad5: q<=8'hb8;
	15'h6ad6: q<=8'h50;
	15'h6ad7: q<=8'h04;
	15'h6ad8: q<=8'ha9;
	15'h6ad9: q<=8'h20;
	15'h6ada: q<=8'h85;
	15'h6adb: q<=8'h4c;
	15'h6adc: q<=8'h20;
	15'h6add: q<=8'h0f;
	15'h6ade: q<=8'hdb;
	15'h6adf: q<=8'h20;
	15'h6ae0: q<=8'h0d;
	15'h6ae1: q<=8'hdf;
	15'h6ae2: q<=8'h8d;
	15'h6ae3: q<=8'h00;
	15'h6ae4: q<=8'h48;
	15'h6ae5: q<=8'he6;
	15'h6ae6: q<=8'h03;
	15'h6ae7: q<=8'ha5;
	15'h6ae8: q<=8'h03;
	15'h6ae9: q<=8'h29;
	15'h6aea: q<=8'h03;
	15'h6aeb: q<=8'hd0;
	15'h6aec: q<=8'h03;
	15'h6aed: q<=8'h20;
	15'h6aee: q<=8'h1b;
	15'h6aef: q<=8'hde;
	15'h6af0: q<=8'had;
	15'h6af1: q<=8'h00;
	15'h6af2: q<=8'h0c;
	15'h6af3: q<=8'h29;
	15'h6af4: q<=8'h10;
	15'h6af5: q<=8'hf0;
	15'h6af6: q<=8'h96;
	15'h6af7: q<=8'hd0;
	15'h6af8: q<=8'hfe;
	15'h6af9: q<=8'h00;
	15'h6afa: q<=8'h04;
	15'h6afb: q<=8'h08;
	15'h6afc: q<=8'h0c;
	15'h6afd: q<=8'h03;
	15'h6afe: q<=8'h07;
	15'h6aff: q<=8'h0b;
	15'h6b00: q<=8'h0b;
	15'h6b01: q<=8'h59;
	15'h6b02: q<=8'hdb;
	15'h6b03: q<=8'hf6;
	15'h6b04: q<=8'hdb;
	15'h6b05: q<=8'h83;
	15'h6b06: q<=8'hdb;
	15'h6b07: q<=8'h99;
	15'h6b08: q<=8'hdb;
	15'h6b09: q<=8'h7d;
	15'h6b0a: q<=8'hdb;
	15'h6b0b: q<=8'h6e;
	15'h6b0c: q<=8'hdb;
	15'h6b0d: q<=8'h21;
	15'h6b0e: q<=8'hdb;
	15'h6b0f: q<=8'ha6;
	15'h6b10: q<=8'h00;
	15'h6b11: q<=8'he0;
	15'h6b12: q<=8'h0e;
	15'h6b13: q<=8'h90;
	15'h6b14: q<=8'h04;
	15'h6b15: q<=8'ha2;
	15'h6b16: q<=8'h02;
	15'h6b17: q<=8'h86;
	15'h6b18: q<=8'h00;
	15'h6b19: q<=8'hbd;
	15'h6b1a: q<=8'h02;
	15'h6b1b: q<=8'hdb;
	15'h6b1c: q<=8'h48;
	15'h6b1d: q<=8'hbd;
	15'h6b1e: q<=8'h01;
	15'h6b1f: q<=8'hdb;
	15'h6b20: q<=8'h48;
	15'h6b21: q<=8'h60;
	15'h6b22: q<=8'ha9;
	15'h6b23: q<=8'h00;
	15'h6b24: q<=8'h8d;
	15'h6b25: q<=8'he0;
	15'h6b26: q<=8'h60;
	15'h6b27: q<=8'h8d;
	15'h6b28: q<=8'h80;
	15'h6b29: q<=8'h60;
	15'h6b2a: q<=8'h8d;
	15'h6b2b: q<=8'hc0;
	15'h6b2c: q<=8'h60;
	15'h6b2d: q<=8'h8d;
	15'h6b2e: q<=8'hd0;
	15'h6b2f: q<=8'h60;
	15'h6b30: q<=8'h8d;
	15'h6b31: q<=8'h00;
	15'h6b32: q<=8'h60;
	15'h6b33: q<=8'h8d;
	15'h6b34: q<=8'h40;
	15'h6b35: q<=8'h60;
	15'h6b36: q<=8'had;
	15'h6b37: q<=8'h40;
	15'h6b38: q<=8'h60;
	15'h6b39: q<=8'had;
	15'h6b3a: q<=8'h60;
	15'h6b3b: q<=8'h60;
	15'h6b3c: q<=8'had;
	15'h6b3d: q<=8'h70;
	15'h6b3e: q<=8'h60;
	15'h6b3f: q<=8'had;
	15'h6b40: q<=8'h50;
	15'h6b41: q<=8'h60;
	15'h6b42: q<=8'ha9;
	15'h6b43: q<=8'h08;
	15'h6b44: q<=8'h8d;
	15'h6b45: q<=8'he0;
	15'h6b46: q<=8'h60;
	15'h6b47: q<=8'ha9;
	15'h6b48: q<=8'h01;
	15'h6b49: q<=8'ha2;
	15'h6b4a: q<=8'h1f;
	15'h6b4b: q<=8'h18;
	15'h6b4c: q<=8'h9d;
	15'h6b4d: q<=8'h80;
	15'h6b4e: q<=8'h60;
	15'h6b4f: q<=8'h2a;
	15'h6b50: q<=8'hca;
	15'h6b51: q<=8'h10;
	15'h6b52: q<=8'hf9;
	15'h6b53: q<=8'ha9;
	15'h6b54: q<=8'h34;
	15'h6b55: q<=8'ha2;
	15'h6b56: q<=8'ha6;
	15'h6b57: q<=8'h4c;
	15'h6b58: q<=8'h39;
	15'h6b59: q<=8'hdf;
	15'h6b5a: q<=8'had;
	15'h6b5b: q<=8'hca;
	15'h6b5c: q<=8'h01;
	15'h6b5d: q<=8'h0d;
	15'h6b5e: q<=8'hc7;
	15'h6b5f: q<=8'h01;
	15'h6b60: q<=8'hd0;
	15'h6b61: q<=8'h0c;
	15'h6b62: q<=8'h20;
	15'h6b63: q<=8'h11;
	15'h6b64: q<=8'hde;
	15'h6b65: q<=8'had;
	15'h6b66: q<=8'hc9;
	15'h6b67: q<=8'h01;
	15'h6b68: q<=8'h85;
	15'h6b69: q<=8'h7c;
	15'h6b6a: q<=8'ha9;
	15'h6b6b: q<=8'h02;
	15'h6b6c: q<=8'h85;
	15'h6b6d: q<=8'h00;
	15'h6b6e: q<=8'h60;
	15'h6b6f: q<=8'ha5;
	15'h6b70: q<=8'h50;
	15'h6b71: q<=8'h4a;
	15'h6b72: q<=8'ha8;
	15'h6b73: q<=8'ha9;
	15'h6b74: q<=8'h68;
	15'h6b75: q<=8'h20;
	15'h6b76: q<=8'h4c;
	15'h6b77: q<=8'hdf;
	15'h6b78: q<=8'ha2;
	15'h6b79: q<=8'h4e;
	15'h6b7a: q<=8'ha9;
	15'h6b7b: q<=8'h33;
	15'h6b7c: q<=8'hd0;
	15'h6b7d: q<=8'h0a;
	15'h6b7e: q<=8'ha2;
	15'h6b7f: q<=8'hb6;
	15'h6b80: q<=8'ha9;
	15'h6b81: q<=8'h32;
	15'h6b82: q<=8'hd0;
	15'h6b83: q<=8'h04;
	15'h6b84: q<=8'ha9;
	15'h6b85: q<=8'h33;
	15'h6b86: q<=8'ha2;
	15'h6b87: q<=8'h0a;
	15'h6b88: q<=8'h20;
	15'h6b89: q<=8'h39;
	15'h6b8a: q<=8'hdf;
	15'h6b8b: q<=8'ha2;
	15'h6b8c: q<=8'h06;
	15'h6b8d: q<=8'ha9;
	15'h6b8e: q<=8'h00;
	15'h6b8f: q<=8'h9d;
	15'h6b90: q<=8'hc1;
	15'h6b91: q<=8'h60;
	15'h6b92: q<=8'h9d;
	15'h6b93: q<=8'hd1;
	15'h6b94: q<=8'h60;
	15'h6b95: q<=8'hca;
	15'h6b96: q<=8'hca;
	15'h6b97: q<=8'h10;
	15'h6b98: q<=8'hf6;
	15'h6b99: q<=8'h60;
	15'h6b9a: q<=8'ha5;
	15'h6b9b: q<=8'h03;
	15'h6b9c: q<=8'h29;
	15'h6b9d: q<=8'h3f;
	15'h6b9e: q<=8'hd0;
	15'h6b9f: q<=8'h02;
	15'h6ba0: q<=8'he6;
	15'h6ba1: q<=8'h39;
	15'h6ba2: q<=8'ha5;
	15'h6ba3: q<=8'h39;
	15'h6ba4: q<=8'h29;
	15'h6ba5: q<=8'h07;
	15'h6ba6: q<=8'haa;
	15'h6ba7: q<=8'hbc;
	15'h6ba8: q<=8'hd5;
	15'h6ba9: q<=8'hdb;
	15'h6baa: q<=8'ha9;
	15'h6bab: q<=8'h00;
	15'h6bac: q<=8'h99;
	15'h6bad: q<=8'hc1;
	15'h6bae: q<=8'h60;
	15'h6baf: q<=8'hbc;
	15'h6bb0: q<=8'hd6;
	15'h6bb1: q<=8'hdb;
	15'h6bb2: q<=8'hbd;
	15'h6bb3: q<=8'hdc;
	15'h6bb4: q<=8'hdf;
	15'h6bb5: q<=8'h99;
	15'h6bb6: q<=8'hc0;
	15'h6bb7: q<=8'h60;
	15'h6bb8: q<=8'ha9;
	15'h6bb9: q<=8'ha8;
	15'h6bba: q<=8'h99;
	15'h6bbb: q<=8'hc1;
	15'h6bbc: q<=8'h60;
	15'h6bbd: q<=8'ha9;
	15'h6bbe: q<=8'h34;
	15'h6bbf: q<=8'ha2;
	15'h6bc0: q<=8'h56;
	15'h6bc1: q<=8'h20;
	15'h6bc2: q<=8'h39;
	15'h6bc3: q<=8'hdf;
	15'h6bc4: q<=8'ha5;
	15'h6bc5: q<=8'h03;
	15'h6bc6: q<=8'h29;
	15'h6bc7: q<=8'h7f;
	15'h6bc8: q<=8'ha8;
	15'h6bc9: q<=8'ha9;
	15'h6bca: q<=8'h01;
	15'h6bcb: q<=8'h20;
	15'h6bcc: q<=8'h6c;
	15'h6bcd: q<=8'hdf;
	15'h6bce: q<=8'ha9;
	15'h6bcf: q<=8'h34;
	15'h6bd0: q<=8'ha2;
	15'h6bd1: q<=8'haa;
	15'h6bd2: q<=8'h4c;
	15'h6bd3: q<=8'h39;
	15'h6bd4: q<=8'hdf;
	15'h6bd5: q<=8'h16;
	15'h6bd6: q<=8'h00;
	15'h6bd7: q<=8'h10;
	15'h6bd8: q<=8'h02;
	15'h6bd9: q<=8'h12;
	15'h6bda: q<=8'h04;
	15'h6bdb: q<=8'h14;
	15'h6bdc: q<=8'h06;
	15'h6bdd: q<=8'h16;
	15'h6bde: q<=8'h00;
	15'h6bdf: q<=8'hea;
	15'h6be0: q<=8'h8d;
	15'h6be1: q<=8'hdb;
	15'h6be2: q<=8'h60;
	15'h6be3: q<=8'had;
	15'h6be4: q<=8'hd8;
	15'h6be5: q<=8'h60;
	15'h6be6: q<=8'h29;
	15'h6be7: q<=8'h07;
	15'h6be8: q<=8'h85;
	15'h6be9: q<=8'h37;
	15'h6bea: q<=8'h8d;
	15'h6beb: q<=8'hcb;
	15'h6bec: q<=8'h60;
	15'h6bed: q<=8'had;
	15'h6bee: q<=8'hc8;
	15'h6bef: q<=8'h60;
	15'h6bf0: q<=8'h29;
	15'h6bf1: q<=8'h20;
	15'h6bf2: q<=8'h4a;
	15'h6bf3: q<=8'h4a;
	15'h6bf4: q<=8'h05;
	15'h6bf5: q<=8'h37;
	15'h6bf6: q<=8'h60;
	15'h6bf7: q<=8'ha5;
	15'h6bf8: q<=8'h2e;
	15'h6bf9: q<=8'hf0;
	15'h6bfa: q<=8'h1e;
	15'h6bfb: q<=8'h8d;
	15'h6bfc: q<=8'h95;
	15'h6bfd: q<=8'h60;
	15'h6bfe: q<=8'h8d;
	15'h6bff: q<=8'h8d;
	15'h6c00: q<=8'h60;
	15'h6c01: q<=8'ha5;
	15'h6c02: q<=8'h2f;
	15'h6c03: q<=8'h8d;
	15'h6c04: q<=8'h96;
	15'h6c05: q<=8'h60;
	15'h6c06: q<=8'ha2;
	15'h6c07: q<=8'h00;
	15'h6c08: q<=8'h20;
	15'h6c09: q<=8'he6;
	15'h6c0a: q<=8'hdc;
	15'h6c0b: q<=8'hc9;
	15'h6c0c: q<=8'h01;
	15'h6c0d: q<=8'hd0;
	15'h6c0e: q<=8'h06;
	15'h6c0f: q<=8'h98;
	15'h6c10: q<=8'hd0;
	15'h6c11: q<=8'h03;
	15'h6c12: q<=8'h8a;
	15'h6c13: q<=8'h10;
	15'h6c14: q<=8'h04;
	15'h6c15: q<=8'ha9;
	15'h6c16: q<=8'hff;
	15'h6c17: q<=8'h85;
	15'h6c18: q<=8'h78;
	15'h6c19: q<=8'ha2;
	15'h6c1a: q<=8'h00;
	15'h6c1b: q<=8'h86;
	15'h6c1c: q<=8'h73;
	15'h6c1d: q<=8'he6;
	15'h6c1e: q<=8'h2e;
	15'h6c1f: q<=8'hd0;
	15'h6c20: q<=8'h06;
	15'h6c21: q<=8'he6;
	15'h6c22: q<=8'h2f;
	15'h6c23: q<=8'h10;
	15'h6c24: q<=8'h02;
	15'h6c25: q<=8'h86;
	15'h6c26: q<=8'h2f;
	15'h6c27: q<=8'h8d;
	15'h6c28: q<=8'hdb;
	15'h6c29: q<=8'h60;
	15'h6c2a: q<=8'had;
	15'h6c2b: q<=8'hd8;
	15'h6c2c: q<=8'h60;
	15'h6c2d: q<=8'h29;
	15'h6c2e: q<=8'h78;
	15'h6c2f: q<=8'h85;
	15'h6c30: q<=8'h4d;
	15'h6c31: q<=8'hf0;
	15'h6c32: q<=8'h05;
	15'h6c33: q<=8'h8d;
	15'h6c34: q<=8'hc0;
	15'h6c35: q<=8'h60;
	15'h6c36: q<=8'ha2;
	15'h6c37: q<=8'ha4;
	15'h6c38: q<=8'h8e;
	15'h6c39: q<=8'hc1;
	15'h6c3a: q<=8'h60;
	15'h6c3b: q<=8'ha2;
	15'h6c3c: q<=8'h00;
	15'h6c3d: q<=8'ha5;
	15'h6c3e: q<=8'h4e;
	15'h6c3f: q<=8'hf0;
	15'h6c40: q<=8'h06;
	15'h6c41: q<=8'h0a;
	15'h6c42: q<=8'h8d;
	15'h6c43: q<=8'hc2;
	15'h6c44: q<=8'h60;
	15'h6c45: q<=8'ha2;
	15'h6c46: q<=8'ha4;
	15'h6c47: q<=8'h8e;
	15'h6c48: q<=8'hc3;
	15'h6c49: q<=8'h60;
	15'h6c4a: q<=8'h20;
	15'h6c4b: q<=8'h0d;
	15'h6c4c: q<=8'hdd;
	15'h6c4d: q<=8'ha4;
	15'h6c4e: q<=8'h4d;
	15'h6c4f: q<=8'ha9;
	15'h6c50: q<=8'hd0;
	15'h6c51: q<=8'ha2;
	15'h6c52: q<=8'hf0;
	15'h6c53: q<=8'h20;
	15'h6c54: q<=8'h2b;
	15'h6c55: q<=8'hdd;
	15'h6c56: q<=8'ha4;
	15'h6c57: q<=8'h4e;
	15'h6c58: q<=8'h20;
	15'h6c59: q<=8'h27;
	15'h6c5a: q<=8'hdd;
	15'h6c5b: q<=8'ha5;
	15'h6c5c: q<=8'h52;
	15'h6c5d: q<=8'h29;
	15'h6c5e: q<=8'h10;
	15'h6c5f: q<=8'hf0;
	15'h6c60: q<=8'h1d;
	15'h6c61: q<=8'ha9;
	15'h6c62: q<=8'h34;
	15'h6c63: q<=8'ha2;
	15'h6c64: q<=8'h82;
	15'h6c65: q<=8'h20;
	15'h6c66: q<=8'h39;
	15'h6c67: q<=8'hdf;
	15'h6c68: q<=8'ha0;
	15'h6c69: q<=8'h10;
	15'h6c6a: q<=8'ha5;
	15'h6c6b: q<=8'h4d;
	15'h6c6c: q<=8'h29;
	15'h6c6d: q<=8'h60;
	15'h6c6e: q<=8'hf0;
	15'h6c6f: q<=8'h0e;
	15'h6c70: q<=8'h49;
	15'h6c71: q<=8'h20;
	15'h6c72: q<=8'hf0;
	15'h6c73: q<=8'h04;
	15'h6c74: q<=8'ha9;
	15'h6c75: q<=8'h04;
	15'h6c76: q<=8'ha0;
	15'h6c77: q<=8'h08;
	15'h6c78: q<=8'h8d;
	15'h6c79: q<=8'he0;
	15'h6c7a: q<=8'h60;
	15'h6c7b: q<=8'h8c;
	15'h6c7c: q<=8'h00;
	15'h6c7d: q<=8'h40;
	15'h6c7e: q<=8'ha9;
	15'h6c7f: q<=8'h34;
	15'h6c80: q<=8'ha2;
	15'h6c81: q<=8'h92;
	15'h6c82: q<=8'h20;
	15'h6c83: q<=8'h39;
	15'h6c84: q<=8'hdf;
	15'h6c85: q<=8'ha2;
	15'h6c86: q<=8'h0b;
	15'h6c87: q<=8'hb5;
	15'h6c88: q<=8'h7d;
	15'h6c89: q<=8'hf0;
	15'h6c8a: q<=8'h19;
	15'h6c8b: q<=8'h85;
	15'h6c8c: q<=8'h35;
	15'h6c8d: q<=8'h86;
	15'h6c8e: q<=8'h38;
	15'h6c8f: q<=8'h8a;
	15'h6c90: q<=8'h20;
	15'h6c91: q<=8'h1f;
	15'h6c92: q<=8'hdf;
	15'h6c93: q<=8'ha0;
	15'h6c94: q<=8'hf4;
	15'h6c95: q<=8'ha2;
	15'h6c96: q<=8'hf4;
	15'h6c97: q<=8'ha5;
	15'h6c98: q<=8'h35;
	15'h6c99: q<=8'h20;
	15'h6c9a: q<=8'ha9;
	15'h6c9b: q<=8'hd8;
	15'h6c9c: q<=8'ha9;
	15'h6c9d: q<=8'h0c;
	15'h6c9e: q<=8'haa;
	15'h6c9f: q<=8'h20;
	15'h6ca0: q<=8'h75;
	15'h6ca1: q<=8'hdf;
	15'h6ca2: q<=8'ha6;
	15'h6ca3: q<=8'h38;
	15'h6ca4: q<=8'hca;
	15'h6ca5: q<=8'h10;
	15'h6ca6: q<=8'he0;
	15'h6ca7: q<=8'h20;
	15'h6ca8: q<=8'h53;
	15'h6ca9: q<=8'hdf;
	15'h6caa: q<=8'ha9;
	15'h6cab: q<=8'h00;
	15'h6cac: q<=8'ha2;
	15'h6cad: q<=8'h16;
	15'h6cae: q<=8'h20;
	15'h6caf: q<=8'h75;
	15'h6cb0: q<=8'hdf;
	15'h6cb1: q<=8'ha2;
	15'h6cb2: q<=8'h04;
	15'h6cb3: q<=8'h86;
	15'h6cb4: q<=8'h37;
	15'h6cb5: q<=8'ha6;
	15'h6cb6: q<=8'h37;
	15'h6cb7: q<=8'ha0;
	15'h6cb8: q<=8'h00;
	15'h6cb9: q<=8'hb5;
	15'h6cba: q<=8'h78;
	15'h6cbb: q<=8'hf0;
	15'h6cbc: q<=8'h03;
	15'h6cbd: q<=8'hbc;
	15'h6cbe: q<=8'he1;
	15'h6cbf: q<=8'hdc;
	15'h6cc0: q<=8'hb9;
	15'h6cc1: q<=8'he4;
	15'h6cc2: q<=8'h31;
	15'h6cc3: q<=8'hbe;
	15'h6cc4: q<=8'he5;
	15'h6cc5: q<=8'h31;
	15'h6cc6: q<=8'h20;
	15'h6cc7: q<=8'h57;
	15'h6cc8: q<=8'hdf;
	15'h6cc9: q<=8'hc6;
	15'h6cca: q<=8'h37;
	15'h6ccb: q<=8'h10;
	15'h6ccc: q<=8'he8;
	15'h6ccd: q<=8'ha2;
	15'h6cce: q<=8'hac;
	15'h6ccf: q<=8'ha9;
	15'h6cd0: q<=8'h30;
	15'h6cd1: q<=8'h20;
	15'h6cd2: q<=8'h75;
	15'h6cd3: q<=8'hdf;
	15'h6cd4: q<=8'ha4;
	15'h6cd5: q<=8'h50;
	15'h6cd6: q<=8'hb9;
	15'h6cd7: q<=8'he8;
	15'h6cd8: q<=8'hdf;
	15'h6cd9: q<=8'hbe;
	15'h6cda: q<=8'he4;
	15'h6cdb: q<=8'hdf;
	15'h6cdc: q<=8'ha0;
	15'h6cdd: q<=8'hc0;
	15'h6cde: q<=8'h4c;
	15'h6cdf: q<=8'h73;
	15'h6ce0: q<=8'hdf;
	15'h6ce1: q<=8'h2e;
	15'h6ce2: q<=8'h38;
	15'h6ce3: q<=8'h34;
	15'h6ce4: q<=8'h36;
	15'h6ce5: q<=8'h1e;
	15'h6ce6: q<=8'ha0;
	15'h6ce7: q<=8'h00;
	15'h6ce8: q<=8'h84;
	15'h6ce9: q<=8'h73;
	15'h6cea: q<=8'h8c;
	15'h6ceb: q<=8'h14;
	15'h6cec: q<=8'h04;
	15'h6ced: q<=8'h8d;
	15'h6cee: q<=8'h8e;
	15'h6cef: q<=8'h60;
	15'h6cf0: q<=8'h8e;
	15'h6cf1: q<=8'h8f;
	15'h6cf2: q<=8'h60;
	15'h6cf3: q<=8'h8c;
	15'h6cf4: q<=8'h90;
	15'h6cf5: q<=8'h60;
	15'h6cf6: q<=8'ha2;
	15'h6cf7: q<=8'h10;
	15'h6cf8: q<=8'h8e;
	15'h6cf9: q<=8'h8c;
	15'h6cfa: q<=8'h60;
	15'h6cfb: q<=8'h8e;
	15'h6cfc: q<=8'h94;
	15'h6cfd: q<=8'h60;
	15'h6cfe: q<=8'hca;
	15'h6cff: q<=8'h30;
	15'h6d00: q<=8'h0b;
	15'h6d01: q<=8'had;
	15'h6d02: q<=8'h40;
	15'h6d03: q<=8'h60;
	15'h6d04: q<=8'h30;
	15'h6d05: q<=8'hf8;
	15'h6d06: q<=8'had;
	15'h6d07: q<=8'h60;
	15'h6d08: q<=8'h60;
	15'h6d09: q<=8'hac;
	15'h6d0a: q<=8'h70;
	15'h6d0b: q<=8'h60;
	15'h6d0c: q<=8'h60;
	15'h6d0d: q<=8'h20;
	15'h6d0e: q<=8'h53;
	15'h6d0f: q<=8'hdf;
	15'h6d10: q<=8'ha9;
	15'h6d11: q<=8'h00;
	15'h6d12: q<=8'h20;
	15'h6d13: q<=8'h6a;
	15'h6d14: q<=8'hdf;
	15'h6d15: q<=8'ha9;
	15'h6d16: q<=8'he8;
	15'h6d17: q<=8'hac;
	15'h6d18: q<=8'h00;
	15'h6d19: q<=8'h0d;
	15'h6d1a: q<=8'h20;
	15'h6d1b: q<=8'h29;
	15'h6d1c: q<=8'hdd;
	15'h6d1d: q<=8'hac;
	15'h6d1e: q<=8'h00;
	15'h6d1f: q<=8'h0e;
	15'h6d20: q<=8'h20;
	15'h6d21: q<=8'h27;
	15'h6d22: q<=8'hdd;
	15'h6d23: q<=8'h20;
	15'h6d24: q<=8'he0;
	15'h6d25: q<=8'hdb;
	15'h6d26: q<=8'ha8;
	15'h6d27: q<=8'ha9;
	15'h6d28: q<=8'hd0;
	15'h6d29: q<=8'ha2;
	15'h6d2a: q<=8'hf8;
	15'h6d2b: q<=8'h84;
	15'h6d2c: q<=8'h35;
	15'h6d2d: q<=8'h20;
	15'h6d2e: q<=8'h75;
	15'h6d2f: q<=8'hdf;
	15'h6d30: q<=8'ha2;
	15'h6d31: q<=8'h07;
	15'h6d32: q<=8'h86;
	15'h6d33: q<=8'h37;
	15'h6d34: q<=8'h06;
	15'h6d35: q<=8'h35;
	15'h6d36: q<=8'ha9;
	15'h6d37: q<=8'h00;
	15'h6d38: q<=8'h2a;
	15'h6d39: q<=8'h20;
	15'h6d3a: q<=8'h1f;
	15'h6d3b: q<=8'hdf;
	15'h6d3c: q<=8'hc6;
	15'h6d3d: q<=8'h37;
	15'h6d3e: q<=8'h10;
	15'h6d3f: q<=8'hf4;
	15'h6d40: q<=8'h60;
	15'h6d41: q<=8'had;
	15'h6d42: q<=8'h0f;
	15'h6d43: q<=8'h04;
	15'h6d44: q<=8'h0a;
	15'h6d45: q<=8'h85;
	15'h6d46: q<=8'h29;
	15'h6d47: q<=8'had;
	15'h6d48: q<=8'h10;
	15'h6d49: q<=8'h04;
	15'h6d4a: q<=8'h2a;
	15'h6d4b: q<=8'h85;
	15'h6d4c: q<=8'h2a;
	15'h6d4d: q<=8'had;
	15'h6d4e: q<=8'h0c;
	15'h6d4f: q<=8'h04;
	15'h6d50: q<=8'h18;
	15'h6d51: q<=8'h65;
	15'h6d52: q<=8'h29;
	15'h6d53: q<=8'h8d;
	15'h6d54: q<=8'h95;
	15'h6d55: q<=8'h60;
	15'h6d56: q<=8'h85;
	15'h6d57: q<=8'h29;
	15'h6d58: q<=8'had;
	15'h6d59: q<=8'h0d;
	15'h6d5a: q<=8'h04;
	15'h6d5b: q<=8'h65;
	15'h6d5c: q<=8'h2a;
	15'h6d5d: q<=8'h8d;
	15'h6d5e: q<=8'h96;
	15'h6d5f: q<=8'h60;
	15'h6d60: q<=8'h05;
	15'h6d61: q<=8'h29;
	15'h6d62: q<=8'hd0;
	15'h6d63: q<=8'h05;
	15'h6d64: q<=8'ha9;
	15'h6d65: q<=8'h01;
	15'h6d66: q<=8'h8d;
	15'h6d67: q<=8'h95;
	15'h6d68: q<=8'h60;
	15'h6d69: q<=8'had;
	15'h6d6a: q<=8'h09;
	15'h6d6b: q<=8'h04;
	15'h6d6c: q<=8'h8d;
	15'h6d6d: q<=8'h8d;
	15'h6d6e: q<=8'h60;
	15'h6d6f: q<=8'had;
	15'h6d70: q<=8'h0a;
	15'h6d71: q<=8'h04;
	15'h6d72: q<=8'hae;
	15'h6d73: q<=8'h0b;
	15'h6d74: q<=8'h04;
	15'h6d75: q<=8'h20;
	15'h6d76: q<=8'he6;
	15'h6d77: q<=8'hdc;
	15'h6d78: q<=8'h8d;
	15'h6d79: q<=8'h12;
	15'h6d7a: q<=8'h04;
	15'h6d7b: q<=8'h8c;
	15'h6d7c: q<=8'h13;
	15'h6d7d: q<=8'h04;
	15'h6d7e: q<=8'ha9;
	15'h6d7f: q<=8'h3d;
	15'h6d80: q<=8'ha2;
	15'h6d81: q<=8'hce;
	15'h6d82: q<=8'h20;
	15'h6d83: q<=8'h39;
	15'h6d84: q<=8'hdf;
	15'h6d85: q<=8'ha9;
	15'h6d86: q<=8'h06;
	15'h6d87: q<=8'h85;
	15'h6d88: q<=8'h3b;
	15'h6d89: q<=8'ha9;
	15'h6d8a: q<=8'h04;
	15'h6d8b: q<=8'h85;
	15'h6d8c: q<=8'h3c;
	15'h6d8d: q<=8'h85;
	15'h6d8e: q<=8'h37;
	15'h6d8f: q<=8'ha0;
	15'h6d90: q<=8'h00;
	15'h6d91: q<=8'h84;
	15'h6d92: q<=8'h31;
	15'h6d93: q<=8'h84;
	15'h6d94: q<=8'h32;
	15'h6d95: q<=8'h84;
	15'h6d96: q<=8'h33;
	15'h6d97: q<=8'h84;
	15'h6d98: q<=8'h34;
	15'h6d99: q<=8'hb1;
	15'h6d9a: q<=8'h3b;
	15'h6d9b: q<=8'h85;
	15'h6d9c: q<=8'h56;
	15'h6d9d: q<=8'he6;
	15'h6d9e: q<=8'h3b;
	15'h6d9f: q<=8'hb1;
	15'h6da0: q<=8'h3b;
	15'h6da1: q<=8'h85;
	15'h6da2: q<=8'h57;
	15'h6da3: q<=8'he6;
	15'h6da4: q<=8'h3b;
	15'h6da5: q<=8'hb1;
	15'h6da6: q<=8'h3b;
	15'h6da7: q<=8'h85;
	15'h6da8: q<=8'h58;
	15'h6da9: q<=8'he6;
	15'h6daa: q<=8'h3b;
	15'h6dab: q<=8'hf8;
	15'h6dac: q<=8'ha0;
	15'h6dad: q<=8'h17;
	15'h6dae: q<=8'h84;
	15'h6daf: q<=8'h38;
	15'h6db0: q<=8'h26;
	15'h6db1: q<=8'h56;
	15'h6db2: q<=8'h26;
	15'h6db3: q<=8'h57;
	15'h6db4: q<=8'h26;
	15'h6db5: q<=8'h58;
	15'h6db6: q<=8'ha0;
	15'h6db7: q<=8'h03;
	15'h6db8: q<=8'ha2;
	15'h6db9: q<=8'h00;
	15'h6dba: q<=8'hb5;
	15'h6dbb: q<=8'h31;
	15'h6dbc: q<=8'h75;
	15'h6dbd: q<=8'h31;
	15'h6dbe: q<=8'h95;
	15'h6dbf: q<=8'h31;
	15'h6dc0: q<=8'he8;
	15'h6dc1: q<=8'h88;
	15'h6dc2: q<=8'h10;
	15'h6dc3: q<=8'hf6;
	15'h6dc4: q<=8'hc6;
	15'h6dc5: q<=8'h38;
	15'h6dc6: q<=8'h10;
	15'h6dc7: q<=8'he8;
	15'h6dc8: q<=8'hd8;
	15'h6dc9: q<=8'ha9;
	15'h6dca: q<=8'h31;
	15'h6dcb: q<=8'ha0;
	15'h6dcc: q<=8'h04;
	15'h6dcd: q<=8'h20;
	15'h6dce: q<=8'hb1;
	15'h6dcf: q<=8'hdf;
	15'h6dd0: q<=8'ha9;
	15'h6dd1: q<=8'hd0;
	15'h6dd2: q<=8'ha2;
	15'h6dd3: q<=8'hf8;
	15'h6dd4: q<=8'h20;
	15'h6dd5: q<=8'h75;
	15'h6dd6: q<=8'hdf;
	15'h6dd7: q<=8'hc6;
	15'h6dd8: q<=8'h37;
	15'h6dd9: q<=8'h10;
	15'h6dda: q<=8'hb4;
	15'h6ddb: q<=8'h60;
	15'h6ddc: q<=8'h73;
	15'h6ddd: q<=8'h00;
	15'h6dde: q<=8'h09;
	15'h6ddf: q<=8'h0a;
	15'h6de0: q<=8'h15;
	15'h6de1: q<=8'h16;
	15'h6de2: q<=8'h22;
	15'h6de3: q<=8'h15;
	15'h6de4: q<=8'h06;
	15'h6de5: q<=8'h15;
	15'h6de6: q<=8'h07;
	15'h6de7: q<=8'h06;
	15'h6de8: q<=8'h04;
	15'h6de9: q<=8'ha9;
	15'h6dea: q<=8'h04;
	15'h6deb: q<=8'hd0;
	15'h6dec: q<=8'h06;
	15'h6ded: q<=8'ha9;
	15'h6dee: q<=8'h03;
	15'h6def: q<=8'hd0;
	15'h6df0: q<=8'h02;
	15'h6df1: q<=8'ha9;
	15'h6df2: q<=8'h07;
	15'h6df3: q<=8'ha0;
	15'h6df4: q<=8'hff;
	15'h6df5: q<=8'hd0;
	15'h6df6: q<=8'h08;
	15'h6df7: q<=8'ha9;
	15'h6df8: q<=8'h03;
	15'h6df9: q<=8'hd0;
	15'h6dfa: q<=8'h02;
	15'h6dfb: q<=8'ha9;
	15'h6dfc: q<=8'h04;
	15'h6dfd: q<=8'ha0;
	15'h6dfe: q<=8'h00;
	15'h6dff: q<=8'h8c;
	15'h6e00: q<=8'hc6;
	15'h6e01: q<=8'h01;
	15'h6e02: q<=8'h48;
	15'h6e03: q<=8'h0d;
	15'h6e04: q<=8'hc7;
	15'h6e05: q<=8'h01;
	15'h6e06: q<=8'h8d;
	15'h6e07: q<=8'hc7;
	15'h6e08: q<=8'h01;
	15'h6e09: q<=8'h68;
	15'h6e0a: q<=8'h0d;
	15'h6e0b: q<=8'hc8;
	15'h6e0c: q<=8'h01;
	15'h6e0d: q<=8'h8d;
	15'h6e0e: q<=8'hc8;
	15'h6e0f: q<=8'h01;
	15'h6e10: q<=8'h60;
	15'h6e11: q<=8'ha9;
	15'h6e12: q<=8'h07;
	15'h6e13: q<=8'h8d;
	15'h6e14: q<=8'hc7;
	15'h6e15: q<=8'h01;
	15'h6e16: q<=8'ha9;
	15'h6e17: q<=8'h00;
	15'h6e18: q<=8'h8d;
	15'h6e19: q<=8'hc8;
	15'h6e1a: q<=8'h01;
	15'h6e1b: q<=8'had;
	15'h6e1c: q<=8'hca;
	15'h6e1d: q<=8'h01;
	15'h6e1e: q<=8'hd0;
	15'h6e1f: q<=8'h4b;
	15'h6e20: q<=8'had;
	15'h6e21: q<=8'hc7;
	15'h6e22: q<=8'h01;
	15'h6e23: q<=8'hf0;
	15'h6e24: q<=8'h46;
	15'h6e25: q<=8'ha2;
	15'h6e26: q<=8'h00;
	15'h6e27: q<=8'h8e;
	15'h6e28: q<=8'hcb;
	15'h6e29: q<=8'h01;
	15'h6e2a: q<=8'h8e;
	15'h6e2b: q<=8'hcf;
	15'h6e2c: q<=8'h01;
	15'h6e2d: q<=8'h8e;
	15'h6e2e: q<=8'hce;
	15'h6e2f: q<=8'h01;
	15'h6e30: q<=8'ha2;
	15'h6e31: q<=8'h08;
	15'h6e32: q<=8'h38;
	15'h6e33: q<=8'h6e;
	15'h6e34: q<=8'hce;
	15'h6e35: q<=8'h01;
	15'h6e36: q<=8'h0a;
	15'h6e37: q<=8'hca;
	15'h6e38: q<=8'h90;
	15'h6e39: q<=8'hf9;
	15'h6e3a: q<=8'ha0;
	15'h6e3b: q<=8'h80;
	15'h6e3c: q<=8'had;
	15'h6e3d: q<=8'hce;
	15'h6e3e: q<=8'h01;
	15'h6e3f: q<=8'h2d;
	15'h6e40: q<=8'hc8;
	15'h6e41: q<=8'h01;
	15'h6e42: q<=8'hd0;
	15'h6e43: q<=8'h02;
	15'h6e44: q<=8'ha0;
	15'h6e45: q<=8'h20;
	15'h6e46: q<=8'h8c;
	15'h6e47: q<=8'hca;
	15'h6e48: q<=8'h01;
	15'h6e49: q<=8'had;
	15'h6e4a: q<=8'hce;
	15'h6e4b: q<=8'h01;
	15'h6e4c: q<=8'h4d;
	15'h6e4d: q<=8'hc7;
	15'h6e4e: q<=8'h01;
	15'h6e4f: q<=8'h8d;
	15'h6e50: q<=8'hc7;
	15'h6e51: q<=8'h01;
	15'h6e52: q<=8'h8a;
	15'h6e53: q<=8'h0a;
	15'h6e54: q<=8'haa;
	15'h6e55: q<=8'hbd;
	15'h6e56: q<=8'hdd;
	15'h6e57: q<=8'hdd;
	15'h6e58: q<=8'h8d;
	15'h6e59: q<=8'hcc;
	15'h6e5a: q<=8'h01;
	15'h6e5b: q<=8'hbd;
	15'h6e5c: q<=8'hde;
	15'h6e5d: q<=8'hdd;
	15'h6e5e: q<=8'h8d;
	15'h6e5f: q<=8'hcd;
	15'h6e60: q<=8'h01;
	15'h6e61: q<=8'hbd;
	15'h6e62: q<=8'he3;
	15'h6e63: q<=8'hdd;
	15'h6e64: q<=8'h85;
	15'h6e65: q<=8'hbd;
	15'h6e66: q<=8'hbd;
	15'h6e67: q<=8'he4;
	15'h6e68: q<=8'hdd;
	15'h6e69: q<=8'h85;
	15'h6e6a: q<=8'hbe;
	15'h6e6b: q<=8'ha0;
	15'h6e6c: q<=8'h00;
	15'h6e6d: q<=8'h8c;
	15'h6e6e: q<=8'h40;
	15'h6e6f: q<=8'h60;
	15'h6e70: q<=8'had;
	15'h6e71: q<=8'hca;
	15'h6e72: q<=8'h01;
	15'h6e73: q<=8'hd0;
	15'h6e74: q<=8'h01;
	15'h6e75: q<=8'h60;
	15'h6e76: q<=8'hac;
	15'h6e77: q<=8'hcb;
	15'h6e78: q<=8'h01;
	15'h6e79: q<=8'hae;
	15'h6e7a: q<=8'hcc;
	15'h6e7b: q<=8'h01;
	15'h6e7c: q<=8'h0a;
	15'h6e7d: q<=8'h90;
	15'h6e7e: q<=8'h0d;
	15'h6e7f: q<=8'h9d;
	15'h6e80: q<=8'h00;
	15'h6e81: q<=8'h60;
	15'h6e82: q<=8'ha9;
	15'h6e83: q<=8'h40;
	15'h6e84: q<=8'h8d;
	15'h6e85: q<=8'hca;
	15'h6e86: q<=8'h01;
	15'h6e87: q<=8'ha0;
	15'h6e88: q<=8'h0e;
	15'h6e89: q<=8'hb8;
	15'h6e8a: q<=8'h50;
	15'h6e8b: q<=8'h73;
	15'h6e8c: q<=8'h10;
	15'h6e8d: q<=8'h25;
	15'h6e8e: q<=8'ha9;
	15'h6e8f: q<=8'h80;
	15'h6e90: q<=8'h8d;
	15'h6e91: q<=8'hca;
	15'h6e92: q<=8'h01;
	15'h6e93: q<=8'had;
	15'h6e94: q<=8'hc6;
	15'h6e95: q<=8'h01;
	15'h6e96: q<=8'hf0;
	15'h6e97: q<=8'h04;
	15'h6e98: q<=8'ha9;
	15'h6e99: q<=8'h00;
	15'h6e9a: q<=8'h91;
	15'h6e9b: q<=8'hbd;
	15'h6e9c: q<=8'hb1;
	15'h6e9d: q<=8'hbd;
	15'h6e9e: q<=8'hec;
	15'h6e9f: q<=8'hcd;
	15'h6ea0: q<=8'h01;
	15'h6ea1: q<=8'h90;
	15'h6ea2: q<=8'h08;
	15'h6ea3: q<=8'ha9;
	15'h6ea4: q<=8'h00;
	15'h6ea5: q<=8'h8d;
	15'h6ea6: q<=8'hca;
	15'h6ea7: q<=8'h01;
	15'h6ea8: q<=8'had;
	15'h6ea9: q<=8'hcf;
	15'h6eaa: q<=8'h01;
	15'h6eab: q<=8'h9d;
	15'h6eac: q<=8'h00;
	15'h6ead: q<=8'h60;
	15'h6eae: q<=8'ha0;
	15'h6eaf: q<=8'h0c;
	15'h6eb0: q<=8'hb8;
	15'h6eb1: q<=8'h50;
	15'h6eb2: q<=8'h3f;
	15'h6eb3: q<=8'ha9;
	15'h6eb4: q<=8'h08;
	15'h6eb5: q<=8'h8d;
	15'h6eb6: q<=8'h40;
	15'h6eb7: q<=8'h60;
	15'h6eb8: q<=8'h9d;
	15'h6eb9: q<=8'h00;
	15'h6eba: q<=8'h60;
	15'h6ebb: q<=8'ha9;
	15'h6ebc: q<=8'h09;
	15'h6ebd: q<=8'h8d;
	15'h6ebe: q<=8'h40;
	15'h6ebf: q<=8'h60;
	15'h6ec0: q<=8'hea;
	15'h6ec1: q<=8'ha9;
	15'h6ec2: q<=8'h08;
	15'h6ec3: q<=8'h8d;
	15'h6ec4: q<=8'h40;
	15'h6ec5: q<=8'h60;
	15'h6ec6: q<=8'hec;
	15'h6ec7: q<=8'hcd;
	15'h6ec8: q<=8'h01;
	15'h6ec9: q<=8'had;
	15'h6eca: q<=8'h50;
	15'h6ecb: q<=8'h60;
	15'h6ecc: q<=8'h90;
	15'h6ecd: q<=8'h20;
	15'h6ece: q<=8'h4d;
	15'h6ecf: q<=8'hcf;
	15'h6ed0: q<=8'h01;
	15'h6ed1: q<=8'hf0;
	15'h6ed2: q<=8'h13;
	15'h6ed3: q<=8'ha9;
	15'h6ed4: q<=8'h00;
	15'h6ed5: q<=8'hac;
	15'h6ed6: q<=8'hcb;
	15'h6ed7: q<=8'h01;
	15'h6ed8: q<=8'h91;
	15'h6ed9: q<=8'hbd;
	15'h6eda: q<=8'h88;
	15'h6edb: q<=8'h10;
	15'h6edc: q<=8'hfb;
	15'h6edd: q<=8'had;
	15'h6ede: q<=8'hce;
	15'h6edf: q<=8'h01;
	15'h6ee0: q<=8'h0d;
	15'h6ee1: q<=8'hc9;
	15'h6ee2: q<=8'h01;
	15'h6ee3: q<=8'h8d;
	15'h6ee4: q<=8'hc9;
	15'h6ee5: q<=8'h01;
	15'h6ee6: q<=8'ha9;
	15'h6ee7: q<=8'h00;
	15'h6ee8: q<=8'h8d;
	15'h6ee9: q<=8'hca;
	15'h6eea: q<=8'h01;
	15'h6eeb: q<=8'hb8;
	15'h6eec: q<=8'h50;
	15'h6eed: q<=8'h02;
	15'h6eee: q<=8'h91;
	15'h6eef: q<=8'hbd;
	15'h6ef0: q<=8'ha0;
	15'h6ef1: q<=8'h00;
	15'h6ef2: q<=8'h18;
	15'h6ef3: q<=8'h6d;
	15'h6ef4: q<=8'hcf;
	15'h6ef5: q<=8'h01;
	15'h6ef6: q<=8'h8d;
	15'h6ef7: q<=8'hcf;
	15'h6ef8: q<=8'h01;
	15'h6ef9: q<=8'hee;
	15'h6efa: q<=8'hcb;
	15'h6efb: q<=8'h01;
	15'h6efc: q<=8'hee;
	15'h6efd: q<=8'hcc;
	15'h6efe: q<=8'h01;
	15'h6eff: q<=8'h8c;
	15'h6f00: q<=8'h40;
	15'h6f01: q<=8'h60;
	15'h6f02: q<=8'h98;
	15'h6f03: q<=8'hd0;
	15'h6f04: q<=8'h03;
	15'h6f05: q<=8'h4c;
	15'h6f06: q<=8'h1b;
	15'h6f07: q<=8'hde;
	15'h6f08: q<=8'h60;
	15'h6f09: q<=8'ha9;
	15'h6f0a: q<=8'hc0;
	15'h6f0b: q<=8'hd0;
	15'h6f0c: q<=8'h05;
	15'h6f0d: q<=8'h20;
	15'h6f0e: q<=8'h53;
	15'h6f0f: q<=8'hdf;
	15'h6f10: q<=8'ha9;
	15'h6f11: q<=8'h20;
	15'h6f12: q<=8'ha0;
	15'h6f13: q<=8'h00;
	15'h6f14: q<=8'h91;
	15'h6f15: q<=8'h74;
	15'h6f16: q<=8'h4c;
	15'h6f17: q<=8'hac;
	15'h6f18: q<=8'hdf;
	15'h6f19: q<=8'h90;
	15'h6f1a: q<=8'h04;
	15'h6f1b: q<=8'h29;
	15'h6f1c: q<=8'h0f;
	15'h6f1d: q<=8'hf0;
	15'h6f1e: q<=8'h05;
	15'h6f1f: q<=8'h29;
	15'h6f20: q<=8'h0f;
	15'h6f21: q<=8'h18;
	15'h6f22: q<=8'h69;
	15'h6f23: q<=8'h01;
	15'h6f24: q<=8'h08;
	15'h6f25: q<=8'h0a;
	15'h6f26: q<=8'ha0;
	15'h6f27: q<=8'h00;
	15'h6f28: q<=8'haa;
	15'h6f29: q<=8'hbd;
	15'h6f2a: q<=8'he4;
	15'h6f2b: q<=8'h31;
	15'h6f2c: q<=8'h91;
	15'h6f2d: q<=8'h74;
	15'h6f2e: q<=8'hbd;
	15'h6f2f: q<=8'he5;
	15'h6f30: q<=8'h31;
	15'h6f31: q<=8'hc8;
	15'h6f32: q<=8'h91;
	15'h6f33: q<=8'h74;
	15'h6f34: q<=8'h20;
	15'h6f35: q<=8'h5f;
	15'h6f36: q<=8'hdf;
	15'h6f37: q<=8'h28;
	15'h6f38: q<=8'h60;
	15'h6f39: q<=8'h4a;
	15'h6f3a: q<=8'h29;
	15'h6f3b: q<=8'h0f;
	15'h6f3c: q<=8'h09;
	15'h6f3d: q<=8'ha0;
	15'h6f3e: q<=8'ha0;
	15'h6f3f: q<=8'h01;
	15'h6f40: q<=8'h91;
	15'h6f41: q<=8'h74;
	15'h6f42: q<=8'h88;
	15'h6f43: q<=8'h8a;
	15'h6f44: q<=8'h6a;
	15'h6f45: q<=8'h91;
	15'h6f46: q<=8'h74;
	15'h6f47: q<=8'hc8;
	15'h6f48: q<=8'hd0;
	15'h6f49: q<=8'h15;
	15'h6f4a: q<=8'ha4;
	15'h6f4b: q<=8'h73;
	15'h6f4c: q<=8'h09;
	15'h6f4d: q<=8'h60;
	15'h6f4e: q<=8'haa;
	15'h6f4f: q<=8'h98;
	15'h6f50: q<=8'h4c;
	15'h6f51: q<=8'h57;
	15'h6f52: q<=8'hdf;
	15'h6f53: q<=8'ha9;
	15'h6f54: q<=8'h40;
	15'h6f55: q<=8'ha2;
	15'h6f56: q<=8'h80;
	15'h6f57: q<=8'ha0;
	15'h6f58: q<=8'h00;
	15'h6f59: q<=8'h91;
	15'h6f5a: q<=8'h74;
	15'h6f5b: q<=8'hc8;
	15'h6f5c: q<=8'h8a;
	15'h6f5d: q<=8'h91;
	15'h6f5e: q<=8'h74;
	15'h6f5f: q<=8'h98;
	15'h6f60: q<=8'h38;
	15'h6f61: q<=8'h65;
	15'h6f62: q<=8'h74;
	15'h6f63: q<=8'h85;
	15'h6f64: q<=8'h74;
	15'h6f65: q<=8'h90;
	15'h6f66: q<=8'h02;
	15'h6f67: q<=8'he6;
	15'h6f68: q<=8'h75;
	15'h6f69: q<=8'h60;
	15'h6f6a: q<=8'ha0;
	15'h6f6b: q<=8'h00;
	15'h6f6c: q<=8'h09;
	15'h6f6d: q<=8'h70;
	15'h6f6e: q<=8'haa;
	15'h6f6f: q<=8'h98;
	15'h6f70: q<=8'h4c;
	15'h6f71: q<=8'h57;
	15'h6f72: q<=8'hdf;
	15'h6f73: q<=8'h84;
	15'h6f74: q<=8'h73;
	15'h6f75: q<=8'ha0;
	15'h6f76: q<=8'h00;
	15'h6f77: q<=8'h0a;
	15'h6f78: q<=8'h90;
	15'h6f79: q<=8'h01;
	15'h6f7a: q<=8'h88;
	15'h6f7b: q<=8'h84;
	15'h6f7c: q<=8'h6f;
	15'h6f7d: q<=8'h0a;
	15'h6f7e: q<=8'h26;
	15'h6f7f: q<=8'h6f;
	15'h6f80: q<=8'h85;
	15'h6f81: q<=8'h6e;
	15'h6f82: q<=8'h8a;
	15'h6f83: q<=8'h0a;
	15'h6f84: q<=8'ha0;
	15'h6f85: q<=8'h00;
	15'h6f86: q<=8'h90;
	15'h6f87: q<=8'h01;
	15'h6f88: q<=8'h88;
	15'h6f89: q<=8'h84;
	15'h6f8a: q<=8'h71;
	15'h6f8b: q<=8'h0a;
	15'h6f8c: q<=8'h26;
	15'h6f8d: q<=8'h71;
	15'h6f8e: q<=8'h85;
	15'h6f8f: q<=8'h70;
	15'h6f90: q<=8'ha2;
	15'h6f91: q<=8'h6e;
	15'h6f92: q<=8'ha0;
	15'h6f93: q<=8'h00;
	15'h6f94: q<=8'hb5;
	15'h6f95: q<=8'h02;
	15'h6f96: q<=8'h91;
	15'h6f97: q<=8'h74;
	15'h6f98: q<=8'hb5;
	15'h6f99: q<=8'h03;
	15'h6f9a: q<=8'h29;
	15'h6f9b: q<=8'h1f;
	15'h6f9c: q<=8'hc8;
	15'h6f9d: q<=8'h91;
	15'h6f9e: q<=8'h74;
	15'h6f9f: q<=8'hb5;
	15'h6fa0: q<=8'h00;
	15'h6fa1: q<=8'hc8;
	15'h6fa2: q<=8'h91;
	15'h6fa3: q<=8'h74;
	15'h6fa4: q<=8'hb5;
	15'h6fa5: q<=8'h01;
	15'h6fa6: q<=8'h45;
	15'h6fa7: q<=8'h73;
	15'h6fa8: q<=8'h29;
	15'h6fa9: q<=8'h1f;
	15'h6faa: q<=8'h45;
	15'h6fab: q<=8'h73;
	15'h6fac: q<=8'hc8;
	15'h6fad: q<=8'h91;
	15'h6fae: q<=8'h74;
	15'h6faf: q<=8'hd0;
	15'h6fb0: q<=8'hae;
	15'h6fb1: q<=8'h38;
	15'h6fb2: q<=8'h08;
	15'h6fb3: q<=8'h88;
	15'h6fb4: q<=8'h84;
	15'h6fb5: q<=8'hae;
	15'h6fb6: q<=8'h18;
	15'h6fb7: q<=8'h65;
	15'h6fb8: q<=8'hae;
	15'h6fb9: q<=8'h28;
	15'h6fba: q<=8'haa;
	15'h6fbb: q<=8'h08;
	15'h6fbc: q<=8'h86;
	15'h6fbd: q<=8'haf;
	15'h6fbe: q<=8'hb5;
	15'h6fbf: q<=8'h00;
	15'h6fc0: q<=8'h4a;
	15'h6fc1: q<=8'h4a;
	15'h6fc2: q<=8'h4a;
	15'h6fc3: q<=8'h4a;
	15'h6fc4: q<=8'h28;
	15'h6fc5: q<=8'h20;
	15'h6fc6: q<=8'h19;
	15'h6fc7: q<=8'hdf;
	15'h6fc8: q<=8'ha5;
	15'h6fc9: q<=8'hae;
	15'h6fca: q<=8'hd0;
	15'h6fcb: q<=8'h01;
	15'h6fcc: q<=8'h18;
	15'h6fcd: q<=8'ha6;
	15'h6fce: q<=8'haf;
	15'h6fcf: q<=8'hb5;
	15'h6fd0: q<=8'h00;
	15'h6fd1: q<=8'h20;
	15'h6fd2: q<=8'h19;
	15'h6fd3: q<=8'hdf;
	15'h6fd4: q<=8'ha6;
	15'h6fd5: q<=8'haf;
	15'h6fd6: q<=8'hca;
	15'h6fd7: q<=8'hc6;
	15'h6fd8: q<=8'hae;
	15'h6fd9: q<=8'h10;
	15'h6fda: q<=8'he0;
	15'h6fdb: q<=8'h60;
	15'h6fdc: q<=8'h10;
	15'h6fdd: q<=8'h10;
	15'h6fde: q<=8'h40;
	15'h6fdf: q<=8'h40;
	15'h6fe0: q<=8'h90;
	15'h6fe1: q<=8'h90;
	15'h6fe2: q<=8'hff;
	15'h6fe3: q<=8'hff;
	15'h6fe4: q<=8'h00;
	15'h6fe5: q<=8'h0c;
	15'h6fe6: q<=8'h16;
	15'h6fe7: q<=8'h1e;
	15'h6fe8: q<=8'h20;
	15'h6fe9: q<=8'h1e;
	15'h6fea: q<=8'h16;
	15'h6feb: q<=8'h0c;
	15'h6fec: q<=8'h00;
	15'h6fed: q<=8'hf4;
	15'h6fee: q<=8'hea;
	15'h6fef: q<=8'he2;
	15'h6ff0: q<=8'he0;
	15'h6ff1: q<=8'he2;
	15'h6ff2: q<=8'hea;
	15'h6ff3: q<=8'hf4;
	15'h6ff4: q<=8'h00;
	15'h6ff5: q<=8'h0c;
	15'h6ff6: q<=8'h16;
	15'h6ff7: q<=8'h1e;
	15'h6ff8: q<=8'h00;
	15'h6ff9: q<=8'h00;
	15'h6ffa: q<=8'h04;
	15'h6ffb: q<=8'hd7;
	15'h6ffc: q<=8'h3f;
	15'h6ffd: q<=8'hd9;
	15'h6ffe: q<=8'h04;
	15'h6fff: q<=8'hd7;
endcase
end
assign dout=q;
endmodule
